magic
tech gf180mcuC
magscale 1 5
timestamp 1670038547
<< obsm1 >>
rect 672 1538 239288 238366
<< metal2 >>
rect 8036 239600 8148 239900
rect 16436 239600 16548 239900
rect 24500 239600 24612 239900
rect 32900 239600 33012 239900
rect 41300 239600 41412 239900
rect 49364 239600 49476 239900
rect 57764 239600 57876 239900
rect 66164 239600 66276 239900
rect 74228 239600 74340 239900
rect 82628 239600 82740 239900
rect 91028 239600 91140 239900
rect 99092 239600 99204 239900
rect 107492 239600 107604 239900
rect 115892 239600 116004 239900
rect 123956 239600 124068 239900
rect 132356 239600 132468 239900
rect 140756 239600 140868 239900
rect 148820 239600 148932 239900
rect 157220 239600 157332 239900
rect 165620 239600 165732 239900
rect 173684 239600 173796 239900
rect 182084 239600 182196 239900
rect 190484 239600 190596 239900
rect 198548 239600 198660 239900
rect 206948 239600 207060 239900
rect 215348 239600 215460 239900
rect 223412 239600 223524 239900
rect 231812 239600 231924 239900
rect 239876 239600 239988 239900
rect -28 100 84 400
rect 8036 100 8148 400
rect 16436 100 16548 400
rect 24500 100 24612 400
rect 32900 100 33012 400
rect 41300 100 41412 400
rect 49364 100 49476 400
rect 57764 100 57876 400
rect 66164 100 66276 400
rect 74228 100 74340 400
rect 82628 100 82740 400
rect 91028 100 91140 400
rect 99092 100 99204 400
rect 107492 100 107604 400
rect 115892 100 116004 400
rect 123956 100 124068 400
rect 132356 100 132468 400
rect 140756 100 140868 400
rect 148820 100 148932 400
rect 157220 100 157332 400
rect 165620 100 165732 400
rect 173684 100 173796 400
rect 182084 100 182196 400
rect 190484 100 190596 400
rect 198548 100 198660 400
rect 206948 100 207060 400
rect 215348 100 215460 400
rect 223412 100 223524 400
rect 231812 100 231924 400
<< obsm2 >>
rect 70 239570 8006 239666
rect 8178 239570 16406 239666
rect 16578 239570 24470 239666
rect 24642 239570 32870 239666
rect 33042 239570 41270 239666
rect 41442 239570 49334 239666
rect 49506 239570 57734 239666
rect 57906 239570 66134 239666
rect 66306 239570 74198 239666
rect 74370 239570 82598 239666
rect 82770 239570 90998 239666
rect 91170 239570 99062 239666
rect 99234 239570 107462 239666
rect 107634 239570 115862 239666
rect 116034 239570 123926 239666
rect 124098 239570 132326 239666
rect 132498 239570 140726 239666
rect 140898 239570 148790 239666
rect 148962 239570 157190 239666
rect 157362 239570 165590 239666
rect 165762 239570 173654 239666
rect 173826 239570 182054 239666
rect 182226 239570 190454 239666
rect 190626 239570 198518 239666
rect 198690 239570 206918 239666
rect 207090 239570 215318 239666
rect 215490 239570 223382 239666
rect 223554 239570 231782 239666
rect 231954 239570 239846 239666
rect 70 430 239890 239570
rect 114 177 8006 430
rect 8178 177 16406 430
rect 16578 177 24470 430
rect 24642 177 32870 430
rect 33042 177 41270 430
rect 41442 177 49334 430
rect 49506 177 57734 430
rect 57906 177 66134 430
rect 66306 177 74198 430
rect 74370 177 82598 430
rect 82770 177 90998 430
rect 91170 177 99062 430
rect 99234 177 107462 430
rect 107634 177 115862 430
rect 116034 177 123926 430
rect 124098 177 132326 430
rect 132498 177 140726 430
rect 140898 177 148790 430
rect 148962 177 157190 430
rect 157362 177 165590 430
rect 165762 177 173654 430
rect 173826 177 182054 430
rect 182226 177 190454 430
rect 190626 177 198518 430
rect 198690 177 206918 430
rect 207090 177 215318 430
rect 215490 177 223382 430
rect 223554 177 231782 430
rect 231954 177 239890 430
<< metal3 >>
rect 100 239876 400 239988
rect 100 231812 400 231924
rect 239600 231812 239900 231924
rect 100 223412 400 223524
rect 239600 223412 239900 223524
rect 100 215348 400 215460
rect 239600 215348 239900 215460
rect 100 206948 400 207060
rect 239600 206948 239900 207060
rect 100 198548 400 198660
rect 239600 198548 239900 198660
rect 100 190484 400 190596
rect 239600 190484 239900 190596
rect 100 182084 400 182196
rect 239600 182084 239900 182196
rect 100 173684 400 173796
rect 239600 173684 239900 173796
rect 100 165620 400 165732
rect 239600 165620 239900 165732
rect 100 157220 400 157332
rect 239600 157220 239900 157332
rect 100 148820 400 148932
rect 239600 148820 239900 148932
rect 100 140756 400 140868
rect 239600 140756 239900 140868
rect 100 132356 400 132468
rect 239600 132356 239900 132468
rect 100 123956 400 124068
rect 239600 123956 239900 124068
rect 100 115892 400 116004
rect 239600 115892 239900 116004
rect 100 107492 400 107604
rect 239600 107492 239900 107604
rect 100 99092 400 99204
rect 239600 99092 239900 99204
rect 100 91028 400 91140
rect 239600 91028 239900 91140
rect 100 82628 400 82740
rect 239600 82628 239900 82740
rect 100 74228 400 74340
rect 239600 74228 239900 74340
rect 100 66164 400 66276
rect 239600 66164 239900 66276
rect 100 57764 400 57876
rect 239600 57764 239900 57876
rect 100 49364 400 49476
rect 239600 49364 239900 49476
rect 100 41300 400 41412
rect 239600 41300 239900 41412
rect 100 32900 400 33012
rect 239600 32900 239900 33012
rect 100 24500 400 24612
rect 239600 24500 239900 24612
rect 100 16436 400 16548
rect 239600 16436 239900 16548
rect 100 8036 400 8148
rect 239600 8036 239900 8148
rect 239600 -28 239900 84
<< obsm3 >>
rect 430 239846 239895 239890
rect 350 231954 239895 239846
rect 430 231782 239570 231954
rect 350 223554 239895 231782
rect 430 223382 239570 223554
rect 350 215490 239895 223382
rect 430 215318 239570 215490
rect 350 207090 239895 215318
rect 430 206918 239570 207090
rect 350 198690 239895 206918
rect 430 198518 239570 198690
rect 350 190626 239895 198518
rect 430 190454 239570 190626
rect 350 182226 239895 190454
rect 430 182054 239570 182226
rect 350 173826 239895 182054
rect 430 173654 239570 173826
rect 350 165762 239895 173654
rect 430 165590 239570 165762
rect 350 157362 239895 165590
rect 430 157190 239570 157362
rect 350 148962 239895 157190
rect 430 148790 239570 148962
rect 350 140898 239895 148790
rect 430 140726 239570 140898
rect 350 132498 239895 140726
rect 430 132326 239570 132498
rect 350 124098 239895 132326
rect 430 123926 239570 124098
rect 350 116034 239895 123926
rect 430 115862 239570 116034
rect 350 107634 239895 115862
rect 430 107462 239570 107634
rect 350 99234 239895 107462
rect 430 99062 239570 99234
rect 350 91170 239895 99062
rect 430 90998 239570 91170
rect 350 82770 239895 90998
rect 430 82598 239570 82770
rect 350 74370 239895 82598
rect 430 74198 239570 74370
rect 350 66306 239895 74198
rect 430 66134 239570 66306
rect 350 57906 239895 66134
rect 430 57734 239570 57906
rect 350 49506 239895 57734
rect 430 49334 239570 49506
rect 350 41442 239895 49334
rect 430 41270 239570 41442
rect 350 33042 239895 41270
rect 430 32870 239570 33042
rect 350 24642 239895 32870
rect 430 24470 239570 24642
rect 350 16578 239895 24470
rect 430 16406 239570 16578
rect 350 8178 239895 16406
rect 430 8006 239570 8178
rect 350 114 239895 8006
rect 350 70 239570 114
<< metal4 >>
rect 2224 1538 2384 238366
rect 9904 1538 10064 238366
rect 17584 1538 17744 238366
rect 25264 1538 25424 238366
rect 32944 1538 33104 238366
rect 40624 1538 40784 238366
rect 48304 1538 48464 238366
rect 55984 1538 56144 238366
rect 63664 1538 63824 238366
rect 71344 1538 71504 238366
rect 79024 1538 79184 238366
rect 86704 1538 86864 238366
rect 94384 1538 94544 238366
rect 102064 1538 102224 238366
rect 109744 1538 109904 238366
rect 117424 1538 117584 238366
rect 125104 1538 125264 238366
rect 132784 1538 132944 238366
rect 140464 1538 140624 238366
rect 148144 1538 148304 238366
rect 155824 1538 155984 238366
rect 163504 1538 163664 238366
rect 171184 1538 171344 238366
rect 178864 1538 179024 238366
rect 186544 1538 186704 238366
rect 194224 1538 194384 238366
rect 201904 1538 202064 238366
rect 209584 1538 209744 238366
rect 217264 1538 217424 238366
rect 224944 1538 225104 238366
rect 232624 1538 232784 238366
<< obsm4 >>
rect 17822 1508 25234 238047
rect 25454 1508 32914 238047
rect 33134 1508 40594 238047
rect 40814 1508 48274 238047
rect 48494 1508 55954 238047
rect 56174 1508 63634 238047
rect 63854 1508 71314 238047
rect 71534 1508 78994 238047
rect 79214 1508 86674 238047
rect 86894 1508 94354 238047
rect 94574 1508 102034 238047
rect 102254 1508 109714 238047
rect 109934 1508 117394 238047
rect 117614 1508 125074 238047
rect 125294 1508 132754 238047
rect 132974 1508 140434 238047
rect 140654 1508 148114 238047
rect 148334 1508 155794 238047
rect 156014 1508 163474 238047
rect 163694 1508 171154 238047
rect 171374 1508 178834 238047
rect 179054 1508 186514 238047
rect 186734 1508 194194 238047
rect 194414 1508 201874 238047
rect 202094 1508 209554 238047
rect 209774 1508 217234 238047
rect 217454 1508 224914 238047
rect 225134 1508 230034 238047
rect 17822 569 230034 1508
<< labels >>
rlabel metal3 s 239600 231812 239900 231924 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 239600 57764 239900 57876 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 24500 239600 24612 239900 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 132356 400 132468 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 215348 239600 215460 239900 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 173684 239600 173796 239900 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 100 148820 400 148932 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 100 41300 400 41412 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 82628 239600 82740 239900 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 66164 100 66276 400 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 100 32900 400 33012 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 239600 215348 239900 215460 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 239600 8036 239900 8148 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 206948 239600 207060 239900 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 100 165620 400 165732 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 100 215348 400 215460 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 239600 107492 239900 107604 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 100 24500 400 24612 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 223412 400 223524 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 115892 239600 116004 239900 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 239600 223412 239900 223524 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 231812 100 231924 400 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 239600 74228 239900 74340 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 107492 239600 107604 239900 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 148820 100 148932 400 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 239600 123956 239900 124068 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 140756 400 140868 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 57764 100 57876 400 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 91028 100 91140 400 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 239600 24500 239900 24612 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 100 182084 400 182196 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 74228 239600 74340 239900 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 239600 82628 239900 82740 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 239600 132356 239900 132468 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 132356 239600 132468 239900 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 239600 99092 239900 99204 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 140756 239600 140868 239900 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 157220 239600 157332 239900 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 190484 239600 190596 239900 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 239876 239600 239988 239900 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 239600 198548 239900 198660 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 32900 100 33012 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 41300 239600 41412 239900 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 107492 100 107604 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 140756 100 140868 400 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 239600 206948 239900 207060 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 215348 100 215460 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 239600 157220 239900 157332 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 99092 239600 99204 239900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 100 115892 400 116004 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 57764 239600 57876 239900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 123956 239600 124068 239900 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 190484 100 190596 400 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 74228 100 74340 400 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 239600 66164 239900 66276 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 66164 239600 66276 239900 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 239600 165620 239900 165732 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 16436 100 16548 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 223412 100 223524 400 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 239600 49364 239900 49476 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 231812 239600 231924 239900 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 100 198548 400 198660 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 198548 100 198660 400 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 99092 100 99204 400 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 100 190484 400 190596 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 239600 182084 239900 182196 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 100 107492 400 107604 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 239600 16436 239900 16548 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 239876 400 239988 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 32900 239600 33012 239900 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 157220 400 157332 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 173684 100 173796 400 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 24500 100 24612 400 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 100 99092 400 99204 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 239600 -28 239900 84 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 239600 140756 239900 140868 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 239600 91028 239900 91140 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 182084 100 182196 400 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 100 173684 400 173796 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 239600 41300 239900 41412 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 123956 400 124068 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 8036 400 8148 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 239600 173684 239900 173796 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 206948 100 207060 400 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 239600 190484 239900 190596 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 123956 100 124068 400 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 100 49364 400 49476 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 100 91028 400 91140 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s -28 100 84 400 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 157220 100 157332 400 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 16436 239600 16548 239900 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 91028 239600 91140 239900 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 165620 239600 165732 239900 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 100 16436 400 16548 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 41300 100 41412 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 8036 100 8148 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 198548 239600 198660 239900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 148820 239600 148932 239900 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 115892 100 116004 400 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 223412 239600 223524 239900 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 239600 32900 239900 33012 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 100 231812 400 231924 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 82628 400 82740 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 49364 100 49476 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 82628 100 82740 400 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 100 74228 400 74340 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 239600 148820 239900 148932 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 132356 100 132468 400 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 100 57764 400 57876 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 182084 239600 182196 239900 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 8036 239600 8148 239900 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 49364 239600 49476 239900 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 165620 100 165732 400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 66164 400 66276 6 io_out[9]
port 114 nsew signal output
rlabel metal4 s 2224 1538 2384 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 238366 6 vdd
port 115 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 238366 6 vss
port 116 nsew ground bidirectional
rlabel metal3 s 100 206948 400 207060 6 wb_clk_i
port 117 nsew signal input
rlabel metal3 s 239600 115892 239900 116004 6 wb_rst_i
port 118 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 240000 240000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 84627874
string GDS_FILE /home/rs2xd/gf180_shuttle/gf180-rc4/openlane/wrapped_rc4/runs/22_12_02_22_12/results/signoff/wrapped_rc4.magic.gds
string GDS_START 509078
<< end >>

