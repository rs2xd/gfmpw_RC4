magic
tech gf180mcuC
magscale 1 5
timestamp 1669818859
<< obsm1 >>
rect 672 855 89320 58561
<< metal2 >>
rect 672 59600 728 60000
rect 1456 59600 1512 60000
rect 2240 59600 2296 60000
rect 3024 59600 3080 60000
rect 3808 59600 3864 60000
rect 4592 59600 4648 60000
rect 5376 59600 5432 60000
rect 6160 59600 6216 60000
rect 6944 59600 7000 60000
rect 7728 59600 7784 60000
rect 8512 59600 8568 60000
rect 9296 59600 9352 60000
rect 10080 59600 10136 60000
rect 10864 59600 10920 60000
rect 11648 59600 11704 60000
rect 12432 59600 12488 60000
rect 13216 59600 13272 60000
rect 14000 59600 14056 60000
rect 14784 59600 14840 60000
rect 15568 59600 15624 60000
rect 16352 59600 16408 60000
rect 17136 59600 17192 60000
rect 17920 59600 17976 60000
rect 18704 59600 18760 60000
rect 19488 59600 19544 60000
rect 20272 59600 20328 60000
rect 21056 59600 21112 60000
rect 21840 59600 21896 60000
rect 22624 59600 22680 60000
rect 23408 59600 23464 60000
rect 24192 59600 24248 60000
rect 24976 59600 25032 60000
rect 25760 59600 25816 60000
rect 26544 59600 26600 60000
rect 27328 59600 27384 60000
rect 28112 59600 28168 60000
rect 28896 59600 28952 60000
rect 29680 59600 29736 60000
rect 30464 59600 30520 60000
rect 31248 59600 31304 60000
rect 32032 59600 32088 60000
rect 32816 59600 32872 60000
rect 33600 59600 33656 60000
rect 34384 59600 34440 60000
rect 35168 59600 35224 60000
rect 35952 59600 36008 60000
rect 36736 59600 36792 60000
rect 37520 59600 37576 60000
rect 38304 59600 38360 60000
rect 39088 59600 39144 60000
rect 39872 59600 39928 60000
rect 40656 59600 40712 60000
rect 41440 59600 41496 60000
rect 42224 59600 42280 60000
rect 43008 59600 43064 60000
rect 43792 59600 43848 60000
rect 44576 59600 44632 60000
rect 45360 59600 45416 60000
rect 46144 59600 46200 60000
rect 46928 59600 46984 60000
rect 47712 59600 47768 60000
rect 48496 59600 48552 60000
rect 49280 59600 49336 60000
rect 50064 59600 50120 60000
rect 50848 59600 50904 60000
rect 51632 59600 51688 60000
rect 52416 59600 52472 60000
rect 53200 59600 53256 60000
rect 53984 59600 54040 60000
rect 54768 59600 54824 60000
rect 55552 59600 55608 60000
rect 56336 59600 56392 60000
rect 57120 59600 57176 60000
rect 57904 59600 57960 60000
rect 58688 59600 58744 60000
rect 59472 59600 59528 60000
rect 60256 59600 60312 60000
rect 61040 59600 61096 60000
rect 61824 59600 61880 60000
rect 62608 59600 62664 60000
rect 63392 59600 63448 60000
rect 64176 59600 64232 60000
rect 64960 59600 65016 60000
rect 65744 59600 65800 60000
rect 66528 59600 66584 60000
rect 67312 59600 67368 60000
rect 68096 59600 68152 60000
rect 68880 59600 68936 60000
rect 69664 59600 69720 60000
rect 70448 59600 70504 60000
rect 71232 59600 71288 60000
rect 72016 59600 72072 60000
rect 72800 59600 72856 60000
rect 73584 59600 73640 60000
rect 74368 59600 74424 60000
rect 75152 59600 75208 60000
rect 75936 59600 75992 60000
rect 76720 59600 76776 60000
rect 77504 59600 77560 60000
rect 78288 59600 78344 60000
rect 79072 59600 79128 60000
rect 79856 59600 79912 60000
rect 80640 59600 80696 60000
rect 81424 59600 81480 60000
rect 82208 59600 82264 60000
rect 82992 59600 83048 60000
rect 83776 59600 83832 60000
rect 84560 59600 84616 60000
rect 85344 59600 85400 60000
rect 86128 59600 86184 60000
rect 86912 59600 86968 60000
rect 87696 59600 87752 60000
rect 88480 59600 88536 60000
rect 89264 59600 89320 60000
rect 2968 0 3024 400
rect 3248 0 3304 400
rect 3528 0 3584 400
rect 3808 0 3864 400
rect 4088 0 4144 400
rect 4368 0 4424 400
rect 4648 0 4704 400
rect 4928 0 4984 400
rect 5208 0 5264 400
rect 5488 0 5544 400
rect 5768 0 5824 400
rect 6048 0 6104 400
rect 6328 0 6384 400
rect 6608 0 6664 400
rect 6888 0 6944 400
rect 7168 0 7224 400
rect 7448 0 7504 400
rect 7728 0 7784 400
rect 8008 0 8064 400
rect 8288 0 8344 400
rect 8568 0 8624 400
rect 8848 0 8904 400
rect 9128 0 9184 400
rect 9408 0 9464 400
rect 9688 0 9744 400
rect 9968 0 10024 400
rect 10248 0 10304 400
rect 10528 0 10584 400
rect 10808 0 10864 400
rect 11088 0 11144 400
rect 11368 0 11424 400
rect 11648 0 11704 400
rect 11928 0 11984 400
rect 12208 0 12264 400
rect 12488 0 12544 400
rect 12768 0 12824 400
rect 13048 0 13104 400
rect 13328 0 13384 400
rect 13608 0 13664 400
rect 13888 0 13944 400
rect 14168 0 14224 400
rect 14448 0 14504 400
rect 14728 0 14784 400
rect 15008 0 15064 400
rect 15288 0 15344 400
rect 15568 0 15624 400
rect 15848 0 15904 400
rect 16128 0 16184 400
rect 16408 0 16464 400
rect 16688 0 16744 400
rect 16968 0 17024 400
rect 17248 0 17304 400
rect 17528 0 17584 400
rect 17808 0 17864 400
rect 18088 0 18144 400
rect 18368 0 18424 400
rect 18648 0 18704 400
rect 18928 0 18984 400
rect 19208 0 19264 400
rect 19488 0 19544 400
rect 19768 0 19824 400
rect 20048 0 20104 400
rect 20328 0 20384 400
rect 20608 0 20664 400
rect 20888 0 20944 400
rect 21168 0 21224 400
rect 21448 0 21504 400
rect 21728 0 21784 400
rect 22008 0 22064 400
rect 22288 0 22344 400
rect 22568 0 22624 400
rect 22848 0 22904 400
rect 23128 0 23184 400
rect 23408 0 23464 400
rect 23688 0 23744 400
rect 23968 0 24024 400
rect 24248 0 24304 400
rect 24528 0 24584 400
rect 24808 0 24864 400
rect 25088 0 25144 400
rect 25368 0 25424 400
rect 25648 0 25704 400
rect 25928 0 25984 400
rect 26208 0 26264 400
rect 26488 0 26544 400
rect 26768 0 26824 400
rect 27048 0 27104 400
rect 27328 0 27384 400
rect 27608 0 27664 400
rect 27888 0 27944 400
rect 28168 0 28224 400
rect 28448 0 28504 400
rect 28728 0 28784 400
rect 29008 0 29064 400
rect 29288 0 29344 400
rect 29568 0 29624 400
rect 29848 0 29904 400
rect 30128 0 30184 400
rect 30408 0 30464 400
rect 30688 0 30744 400
rect 30968 0 31024 400
rect 31248 0 31304 400
rect 31528 0 31584 400
rect 31808 0 31864 400
rect 32088 0 32144 400
rect 32368 0 32424 400
rect 32648 0 32704 400
rect 32928 0 32984 400
rect 33208 0 33264 400
rect 33488 0 33544 400
rect 33768 0 33824 400
rect 34048 0 34104 400
rect 34328 0 34384 400
rect 34608 0 34664 400
rect 34888 0 34944 400
rect 35168 0 35224 400
rect 35448 0 35504 400
rect 35728 0 35784 400
rect 36008 0 36064 400
rect 36288 0 36344 400
rect 36568 0 36624 400
rect 36848 0 36904 400
rect 37128 0 37184 400
rect 37408 0 37464 400
rect 37688 0 37744 400
rect 37968 0 38024 400
rect 38248 0 38304 400
rect 38528 0 38584 400
rect 38808 0 38864 400
rect 39088 0 39144 400
rect 39368 0 39424 400
rect 39648 0 39704 400
rect 39928 0 39984 400
rect 40208 0 40264 400
rect 40488 0 40544 400
rect 40768 0 40824 400
rect 41048 0 41104 400
rect 41328 0 41384 400
rect 41608 0 41664 400
rect 41888 0 41944 400
rect 42168 0 42224 400
rect 42448 0 42504 400
rect 42728 0 42784 400
rect 43008 0 43064 400
rect 43288 0 43344 400
rect 43568 0 43624 400
rect 43848 0 43904 400
rect 44128 0 44184 400
rect 44408 0 44464 400
rect 44688 0 44744 400
rect 44968 0 45024 400
rect 45248 0 45304 400
rect 45528 0 45584 400
rect 45808 0 45864 400
rect 46088 0 46144 400
rect 46368 0 46424 400
rect 46648 0 46704 400
rect 46928 0 46984 400
rect 47208 0 47264 400
rect 47488 0 47544 400
rect 47768 0 47824 400
rect 48048 0 48104 400
rect 48328 0 48384 400
rect 48608 0 48664 400
rect 48888 0 48944 400
rect 49168 0 49224 400
rect 49448 0 49504 400
rect 49728 0 49784 400
rect 50008 0 50064 400
rect 50288 0 50344 400
rect 50568 0 50624 400
rect 50848 0 50904 400
rect 51128 0 51184 400
rect 51408 0 51464 400
rect 51688 0 51744 400
rect 51968 0 52024 400
rect 52248 0 52304 400
rect 52528 0 52584 400
rect 52808 0 52864 400
rect 53088 0 53144 400
rect 53368 0 53424 400
rect 53648 0 53704 400
rect 53928 0 53984 400
rect 54208 0 54264 400
rect 54488 0 54544 400
rect 54768 0 54824 400
rect 55048 0 55104 400
rect 55328 0 55384 400
rect 55608 0 55664 400
rect 55888 0 55944 400
rect 56168 0 56224 400
rect 56448 0 56504 400
rect 56728 0 56784 400
rect 57008 0 57064 400
rect 57288 0 57344 400
rect 57568 0 57624 400
rect 57848 0 57904 400
rect 58128 0 58184 400
rect 58408 0 58464 400
rect 58688 0 58744 400
rect 58968 0 59024 400
rect 59248 0 59304 400
rect 59528 0 59584 400
rect 59808 0 59864 400
rect 60088 0 60144 400
rect 60368 0 60424 400
rect 60648 0 60704 400
rect 60928 0 60984 400
rect 61208 0 61264 400
rect 61488 0 61544 400
rect 61768 0 61824 400
rect 62048 0 62104 400
rect 62328 0 62384 400
rect 62608 0 62664 400
rect 62888 0 62944 400
rect 63168 0 63224 400
rect 63448 0 63504 400
rect 63728 0 63784 400
rect 64008 0 64064 400
rect 64288 0 64344 400
rect 64568 0 64624 400
rect 64848 0 64904 400
rect 65128 0 65184 400
rect 65408 0 65464 400
rect 65688 0 65744 400
rect 65968 0 66024 400
rect 66248 0 66304 400
rect 66528 0 66584 400
rect 66808 0 66864 400
rect 67088 0 67144 400
rect 67368 0 67424 400
rect 67648 0 67704 400
rect 67928 0 67984 400
rect 68208 0 68264 400
rect 68488 0 68544 400
rect 68768 0 68824 400
rect 69048 0 69104 400
rect 69328 0 69384 400
rect 69608 0 69664 400
rect 69888 0 69944 400
rect 70168 0 70224 400
rect 70448 0 70504 400
rect 70728 0 70784 400
rect 71008 0 71064 400
rect 71288 0 71344 400
rect 71568 0 71624 400
rect 71848 0 71904 400
rect 72128 0 72184 400
rect 72408 0 72464 400
rect 72688 0 72744 400
rect 72968 0 73024 400
rect 73248 0 73304 400
rect 73528 0 73584 400
rect 73808 0 73864 400
rect 74088 0 74144 400
rect 74368 0 74424 400
rect 74648 0 74704 400
rect 74928 0 74984 400
rect 75208 0 75264 400
rect 75488 0 75544 400
rect 75768 0 75824 400
rect 76048 0 76104 400
rect 76328 0 76384 400
rect 76608 0 76664 400
rect 76888 0 76944 400
rect 77168 0 77224 400
rect 77448 0 77504 400
rect 77728 0 77784 400
rect 78008 0 78064 400
rect 78288 0 78344 400
rect 78568 0 78624 400
rect 78848 0 78904 400
rect 79128 0 79184 400
rect 79408 0 79464 400
rect 79688 0 79744 400
rect 79968 0 80024 400
rect 80248 0 80304 400
rect 80528 0 80584 400
rect 80808 0 80864 400
rect 81088 0 81144 400
rect 81368 0 81424 400
rect 81648 0 81704 400
rect 81928 0 81984 400
rect 82208 0 82264 400
rect 82488 0 82544 400
rect 82768 0 82824 400
rect 83048 0 83104 400
rect 83328 0 83384 400
rect 83608 0 83664 400
rect 83888 0 83944 400
rect 84168 0 84224 400
rect 84448 0 84504 400
rect 84728 0 84784 400
rect 85008 0 85064 400
rect 85288 0 85344 400
rect 85568 0 85624 400
rect 85848 0 85904 400
rect 86128 0 86184 400
rect 86408 0 86464 400
rect 86688 0 86744 400
rect 86968 0 87024 400
<< obsm2 >>
rect 1542 59570 2210 59600
rect 2326 59570 2994 59600
rect 3110 59570 3778 59600
rect 3894 59570 4562 59600
rect 4678 59570 5346 59600
rect 5462 59570 6130 59600
rect 6246 59570 6914 59600
rect 7030 59570 7698 59600
rect 7814 59570 8482 59600
rect 8598 59570 9266 59600
rect 9382 59570 10050 59600
rect 10166 59570 10834 59600
rect 10950 59570 11618 59600
rect 11734 59570 12402 59600
rect 12518 59570 13186 59600
rect 13302 59570 13970 59600
rect 14086 59570 14754 59600
rect 14870 59570 15538 59600
rect 15654 59570 16322 59600
rect 16438 59570 17106 59600
rect 17222 59570 17890 59600
rect 18006 59570 18674 59600
rect 18790 59570 19458 59600
rect 19574 59570 20242 59600
rect 20358 59570 21026 59600
rect 21142 59570 21810 59600
rect 21926 59570 22594 59600
rect 22710 59570 23378 59600
rect 23494 59570 24162 59600
rect 24278 59570 24946 59600
rect 25062 59570 25730 59600
rect 25846 59570 26514 59600
rect 26630 59570 27298 59600
rect 27414 59570 28082 59600
rect 28198 59570 28866 59600
rect 28982 59570 29650 59600
rect 29766 59570 30434 59600
rect 30550 59570 31218 59600
rect 31334 59570 32002 59600
rect 32118 59570 32786 59600
rect 32902 59570 33570 59600
rect 33686 59570 34354 59600
rect 34470 59570 35138 59600
rect 35254 59570 35922 59600
rect 36038 59570 36706 59600
rect 36822 59570 37490 59600
rect 37606 59570 38274 59600
rect 38390 59570 39058 59600
rect 39174 59570 39842 59600
rect 39958 59570 40626 59600
rect 40742 59570 41410 59600
rect 41526 59570 42194 59600
rect 42310 59570 42978 59600
rect 43094 59570 43762 59600
rect 43878 59570 44546 59600
rect 44662 59570 45330 59600
rect 45446 59570 46114 59600
rect 46230 59570 46898 59600
rect 47014 59570 47682 59600
rect 47798 59570 48466 59600
rect 48582 59570 49250 59600
rect 49366 59570 50034 59600
rect 50150 59570 50818 59600
rect 50934 59570 51602 59600
rect 51718 59570 52386 59600
rect 52502 59570 53170 59600
rect 53286 59570 53954 59600
rect 54070 59570 54738 59600
rect 54854 59570 55522 59600
rect 55638 59570 56306 59600
rect 56422 59570 57090 59600
rect 57206 59570 57874 59600
rect 57990 59570 58658 59600
rect 58774 59570 59442 59600
rect 59558 59570 60226 59600
rect 60342 59570 61010 59600
rect 61126 59570 61794 59600
rect 61910 59570 62578 59600
rect 62694 59570 63362 59600
rect 63478 59570 64146 59600
rect 64262 59570 64930 59600
rect 65046 59570 65714 59600
rect 65830 59570 66498 59600
rect 66614 59570 67282 59600
rect 67398 59570 68066 59600
rect 68182 59570 68850 59600
rect 68966 59570 69634 59600
rect 69750 59570 70418 59600
rect 70534 59570 71202 59600
rect 71318 59570 71986 59600
rect 72102 59570 72770 59600
rect 72886 59570 73554 59600
rect 73670 59570 74338 59600
rect 74454 59570 75122 59600
rect 75238 59570 75906 59600
rect 76022 59570 76690 59600
rect 76806 59570 77474 59600
rect 77590 59570 78258 59600
rect 78374 59570 79042 59600
rect 79158 59570 79826 59600
rect 79942 59570 80610 59600
rect 80726 59570 81394 59600
rect 81510 59570 82178 59600
rect 82294 59570 82962 59600
rect 83078 59570 83746 59600
rect 83862 59570 84530 59600
rect 84646 59570 85314 59600
rect 85430 59570 86098 59600
rect 86214 59570 86882 59600
rect 86998 59570 87666 59600
rect 87782 59570 88450 59600
rect 88566 59570 89234 59600
rect 1470 430 89306 59570
rect 1470 345 2938 430
rect 3054 345 3218 430
rect 3334 345 3498 430
rect 3614 345 3778 430
rect 3894 345 4058 430
rect 4174 345 4338 430
rect 4454 345 4618 430
rect 4734 345 4898 430
rect 5014 345 5178 430
rect 5294 345 5458 430
rect 5574 345 5738 430
rect 5854 345 6018 430
rect 6134 345 6298 430
rect 6414 345 6578 430
rect 6694 345 6858 430
rect 6974 345 7138 430
rect 7254 345 7418 430
rect 7534 345 7698 430
rect 7814 345 7978 430
rect 8094 345 8258 430
rect 8374 345 8538 430
rect 8654 345 8818 430
rect 8934 345 9098 430
rect 9214 345 9378 430
rect 9494 345 9658 430
rect 9774 345 9938 430
rect 10054 345 10218 430
rect 10334 345 10498 430
rect 10614 345 10778 430
rect 10894 345 11058 430
rect 11174 345 11338 430
rect 11454 345 11618 430
rect 11734 345 11898 430
rect 12014 345 12178 430
rect 12294 345 12458 430
rect 12574 345 12738 430
rect 12854 345 13018 430
rect 13134 345 13298 430
rect 13414 345 13578 430
rect 13694 345 13858 430
rect 13974 345 14138 430
rect 14254 345 14418 430
rect 14534 345 14698 430
rect 14814 345 14978 430
rect 15094 345 15258 430
rect 15374 345 15538 430
rect 15654 345 15818 430
rect 15934 345 16098 430
rect 16214 345 16378 430
rect 16494 345 16658 430
rect 16774 345 16938 430
rect 17054 345 17218 430
rect 17334 345 17498 430
rect 17614 345 17778 430
rect 17894 345 18058 430
rect 18174 345 18338 430
rect 18454 345 18618 430
rect 18734 345 18898 430
rect 19014 345 19178 430
rect 19294 345 19458 430
rect 19574 345 19738 430
rect 19854 345 20018 430
rect 20134 345 20298 430
rect 20414 345 20578 430
rect 20694 345 20858 430
rect 20974 345 21138 430
rect 21254 345 21418 430
rect 21534 345 21698 430
rect 21814 345 21978 430
rect 22094 345 22258 430
rect 22374 345 22538 430
rect 22654 345 22818 430
rect 22934 345 23098 430
rect 23214 345 23378 430
rect 23494 345 23658 430
rect 23774 345 23938 430
rect 24054 345 24218 430
rect 24334 345 24498 430
rect 24614 345 24778 430
rect 24894 345 25058 430
rect 25174 345 25338 430
rect 25454 345 25618 430
rect 25734 345 25898 430
rect 26014 345 26178 430
rect 26294 345 26458 430
rect 26574 345 26738 430
rect 26854 345 27018 430
rect 27134 345 27298 430
rect 27414 345 27578 430
rect 27694 345 27858 430
rect 27974 345 28138 430
rect 28254 345 28418 430
rect 28534 345 28698 430
rect 28814 345 28978 430
rect 29094 345 29258 430
rect 29374 345 29538 430
rect 29654 345 29818 430
rect 29934 345 30098 430
rect 30214 345 30378 430
rect 30494 345 30658 430
rect 30774 345 30938 430
rect 31054 345 31218 430
rect 31334 345 31498 430
rect 31614 345 31778 430
rect 31894 345 32058 430
rect 32174 345 32338 430
rect 32454 345 32618 430
rect 32734 345 32898 430
rect 33014 345 33178 430
rect 33294 345 33458 430
rect 33574 345 33738 430
rect 33854 345 34018 430
rect 34134 345 34298 430
rect 34414 345 34578 430
rect 34694 345 34858 430
rect 34974 345 35138 430
rect 35254 345 35418 430
rect 35534 345 35698 430
rect 35814 345 35978 430
rect 36094 345 36258 430
rect 36374 345 36538 430
rect 36654 345 36818 430
rect 36934 345 37098 430
rect 37214 345 37378 430
rect 37494 345 37658 430
rect 37774 345 37938 430
rect 38054 345 38218 430
rect 38334 345 38498 430
rect 38614 345 38778 430
rect 38894 345 39058 430
rect 39174 345 39338 430
rect 39454 345 39618 430
rect 39734 345 39898 430
rect 40014 345 40178 430
rect 40294 345 40458 430
rect 40574 345 40738 430
rect 40854 345 41018 430
rect 41134 345 41298 430
rect 41414 345 41578 430
rect 41694 345 41858 430
rect 41974 345 42138 430
rect 42254 345 42418 430
rect 42534 345 42698 430
rect 42814 345 42978 430
rect 43094 345 43258 430
rect 43374 345 43538 430
rect 43654 345 43818 430
rect 43934 345 44098 430
rect 44214 345 44378 430
rect 44494 345 44658 430
rect 44774 345 44938 430
rect 45054 345 45218 430
rect 45334 345 45498 430
rect 45614 345 45778 430
rect 45894 345 46058 430
rect 46174 345 46338 430
rect 46454 345 46618 430
rect 46734 345 46898 430
rect 47014 345 47178 430
rect 47294 345 47458 430
rect 47574 345 47738 430
rect 47854 345 48018 430
rect 48134 345 48298 430
rect 48414 345 48578 430
rect 48694 345 48858 430
rect 48974 345 49138 430
rect 49254 345 49418 430
rect 49534 345 49698 430
rect 49814 345 49978 430
rect 50094 345 50258 430
rect 50374 345 50538 430
rect 50654 345 50818 430
rect 50934 345 51098 430
rect 51214 345 51378 430
rect 51494 345 51658 430
rect 51774 345 51938 430
rect 52054 345 52218 430
rect 52334 345 52498 430
rect 52614 345 52778 430
rect 52894 345 53058 430
rect 53174 345 53338 430
rect 53454 345 53618 430
rect 53734 345 53898 430
rect 54014 345 54178 430
rect 54294 345 54458 430
rect 54574 345 54738 430
rect 54854 345 55018 430
rect 55134 345 55298 430
rect 55414 345 55578 430
rect 55694 345 55858 430
rect 55974 345 56138 430
rect 56254 345 56418 430
rect 56534 345 56698 430
rect 56814 345 56978 430
rect 57094 345 57258 430
rect 57374 345 57538 430
rect 57654 345 57818 430
rect 57934 345 58098 430
rect 58214 345 58378 430
rect 58494 345 58658 430
rect 58774 345 58938 430
rect 59054 345 59218 430
rect 59334 345 59498 430
rect 59614 345 59778 430
rect 59894 345 60058 430
rect 60174 345 60338 430
rect 60454 345 60618 430
rect 60734 345 60898 430
rect 61014 345 61178 430
rect 61294 345 61458 430
rect 61574 345 61738 430
rect 61854 345 62018 430
rect 62134 345 62298 430
rect 62414 345 62578 430
rect 62694 345 62858 430
rect 62974 345 63138 430
rect 63254 345 63418 430
rect 63534 345 63698 430
rect 63814 345 63978 430
rect 64094 345 64258 430
rect 64374 345 64538 430
rect 64654 345 64818 430
rect 64934 345 65098 430
rect 65214 345 65378 430
rect 65494 345 65658 430
rect 65774 345 65938 430
rect 66054 345 66218 430
rect 66334 345 66498 430
rect 66614 345 66778 430
rect 66894 345 67058 430
rect 67174 345 67338 430
rect 67454 345 67618 430
rect 67734 345 67898 430
rect 68014 345 68178 430
rect 68294 345 68458 430
rect 68574 345 68738 430
rect 68854 345 69018 430
rect 69134 345 69298 430
rect 69414 345 69578 430
rect 69694 345 69858 430
rect 69974 345 70138 430
rect 70254 345 70418 430
rect 70534 345 70698 430
rect 70814 345 70978 430
rect 71094 345 71258 430
rect 71374 345 71538 430
rect 71654 345 71818 430
rect 71934 345 72098 430
rect 72214 345 72378 430
rect 72494 345 72658 430
rect 72774 345 72938 430
rect 73054 345 73218 430
rect 73334 345 73498 430
rect 73614 345 73778 430
rect 73894 345 74058 430
rect 74174 345 74338 430
rect 74454 345 74618 430
rect 74734 345 74898 430
rect 75014 345 75178 430
rect 75294 345 75458 430
rect 75574 345 75738 430
rect 75854 345 76018 430
rect 76134 345 76298 430
rect 76414 345 76578 430
rect 76694 345 76858 430
rect 76974 345 77138 430
rect 77254 345 77418 430
rect 77534 345 77698 430
rect 77814 345 77978 430
rect 78094 345 78258 430
rect 78374 345 78538 430
rect 78654 345 78818 430
rect 78934 345 79098 430
rect 79214 345 79378 430
rect 79494 345 79658 430
rect 79774 345 79938 430
rect 80054 345 80218 430
rect 80334 345 80498 430
rect 80614 345 80778 430
rect 80894 345 81058 430
rect 81174 345 81338 430
rect 81454 345 81618 430
rect 81734 345 81898 430
rect 82014 345 82178 430
rect 82294 345 82458 430
rect 82574 345 82738 430
rect 82854 345 83018 430
rect 83134 345 83298 430
rect 83414 345 83578 430
rect 83694 345 83858 430
rect 83974 345 84138 430
rect 84254 345 84418 430
rect 84534 345 84698 430
rect 84814 345 84978 430
rect 85094 345 85258 430
rect 85374 345 85538 430
rect 85654 345 85818 430
rect 85934 345 86098 430
rect 86214 345 86378 430
rect 86494 345 86658 430
rect 86774 345 86938 430
rect 87054 345 89306 430
<< obsm3 >>
rect 1465 350 89311 58618
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 28574 1508 32914 58119
rect 33134 1508 40594 58119
rect 40814 1508 48274 58119
rect 48494 1508 55954 58119
rect 56174 1508 63634 58119
rect 63854 1508 70266 58119
rect 28574 1465 70266 1508
<< labels >>
rlabel metal2 s 672 59600 728 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24192 59600 24248 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26544 59600 26600 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28896 59600 28952 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31248 59600 31304 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33600 59600 33656 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 35952 59600 36008 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38304 59600 38360 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40656 59600 40712 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43008 59600 43064 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45360 59600 45416 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3024 59600 3080 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 59600 47768 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52416 59600 52472 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54768 59600 54824 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57120 59600 57176 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 59472 59600 59528 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 61824 59600 61880 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64176 59600 64232 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 66528 59600 66584 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 68880 59600 68936 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5376 59600 5432 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71232 59600 71288 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 73584 59600 73640 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 75936 59600 75992 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 78288 59600 78344 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 80640 59600 80696 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 82992 59600 83048 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 85344 59600 85400 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 87696 59600 87752 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7728 59600 7784 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10080 59600 10136 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12432 59600 12488 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14784 59600 14840 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17136 59600 17192 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19488 59600 19544 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21840 59600 21896 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1456 59600 1512 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 24976 59600 25032 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27328 59600 27384 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32032 59600 32088 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36736 59600 36792 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39088 59600 39144 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41440 59600 41496 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43792 59600 43848 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46144 59600 46200 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3808 59600 3864 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48496 59600 48552 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50848 59600 50904 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53200 59600 53256 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 55552 59600 55608 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57904 59600 57960 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60256 59600 60312 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62608 59600 62664 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 64960 59600 65016 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 67312 59600 67368 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 69664 59600 69720 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6160 59600 6216 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72016 59600 72072 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 74368 59600 74424 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 76720 59600 76776 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79072 59600 79128 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 81424 59600 81480 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 83776 59600 83832 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 86128 59600 86184 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 88480 59600 88536 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8512 59600 8568 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10864 59600 10920 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13216 59600 13272 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17920 59600 17976 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20272 59600 20328 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22624 59600 22680 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2240 59600 2296 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25760 59600 25816 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28112 59600 28168 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30464 59600 30520 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32816 59600 32872 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35168 59600 35224 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 39872 59600 39928 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42224 59600 42280 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46928 59600 46984 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4592 59600 4648 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49280 59600 49336 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51632 59600 51688 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53984 59600 54040 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56336 59600 56392 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61040 59600 61096 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63392 59600 63448 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 65744 59600 65800 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68096 59600 68152 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 70448 59600 70504 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6944 59600 7000 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 72800 59600 72856 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75152 59600 75208 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 77504 59600 77560 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 79856 59600 79912 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 82208 59600 82264 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 84560 59600 84616 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 86912 59600 86968 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 89264 59600 89320 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11648 59600 11704 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14000 59600 14056 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18704 59600 18760 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21056 59600 21112 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86408 0 86464 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 86688 0 86744 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 86968 0 87024 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 32648 0 32704 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 41048 0 41104 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 42728 0 42784 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 44408 0 44464 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 46088 0 46144 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 47768 0 47824 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 49448 0 49504 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 51128 0 51184 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 51968 0 52024 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 52808 0 52864 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 54488 0 54544 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 56168 0 56224 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 34328 0 34384 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 57848 0 57904 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 58688 0 58744 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 59528 0 59584 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 61208 0 61264 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 62888 0 62944 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 64568 0 64624 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 65408 0 65464 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 66248 0 66304 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 67088 0 67144 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 67928 0 67984 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 68768 0 68824 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 69608 0 69664 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 70448 0 70504 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 71288 0 71344 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 72968 0 73024 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 73808 0 73864 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 36008 0 36064 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 74648 0 74704 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 76328 0 76384 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 78008 0 78064 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 78848 0 78904 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 79688 0 79744 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 80528 0 80584 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 81368 0 81424 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 82208 0 82264 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 83048 0 83104 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 84728 0 84784 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 85568 0 85624 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 37688 0 37744 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 39368 0 39424 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 42168 0 42224 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 43008 0 43064 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 43848 0 43904 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 44688 0 44744 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 45528 0 45584 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 47208 0 47264 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 48888 0 48944 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 33768 0 33824 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 49728 0 49784 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 50568 0 50624 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 51408 0 51464 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 52248 0 52304 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 53928 0 53984 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 55608 0 55664 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 57288 0 57344 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 58128 0 58184 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 58968 0 59024 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 60648 0 60704 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 62328 0 62384 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 64008 0 64064 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 64848 0 64904 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 65688 0 65744 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 35448 0 35504 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 66528 0 66584 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 67368 0 67424 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 68208 0 68264 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 69048 0 69104 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 69888 0 69944 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 70728 0 70784 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 71568 0 71624 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 72408 0 72464 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 73248 0 73304 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 74088 0 74144 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 74928 0 74984 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 75768 0 75824 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 76608 0 76664 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 77448 0 77504 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 78288 0 78344 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 79128 0 79184 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 79968 0 80024 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 80808 0 80864 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 81648 0 81704 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 82488 0 82544 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 37128 0 37184 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 83328 0 83384 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 84168 0 84224 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 85848 0 85904 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 37968 0 38024 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 38808 0 38864 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 39648 0 39704 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 40488 0 40544 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 33208 0 33264 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 41608 0 41664 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 43288 0 43344 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 46648 0 46704 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 48328 0 48384 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 51688 0 51744 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 53368 0 53424 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 55048 0 55104 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 55888 0 55944 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 56728 0 56784 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 58408 0 58464 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 60088 0 60144 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 60928 0 60984 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 61768 0 61824 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 62608 0 62664 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 63448 0 63504 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 65128 0 65184 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 66808 0 66864 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 68488 0 68544 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 70168 0 70224 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 71848 0 71904 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 73528 0 73584 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 36568 0 36624 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 75208 0 75264 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 76048 0 76104 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 76888 0 76944 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 78568 0 78624 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 80248 0 80304 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 81928 0 81984 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 82768 0 82824 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 83608 0 83664 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 38248 0 38304 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal2 s 2968 0 3024 400 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 3248 0 3304 400 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 3528 0 3584 400 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 4648 0 4704 400 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 14168 0 14224 400 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 15848 0 15904 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 17528 0 17584 400 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 19208 0 19264 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 20888 0 20944 400 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 5768 0 5824 400 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 22568 0 22624 400 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 24248 0 24304 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 25928 0 25984 400 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 27608 0 27664 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 29288 0 29344 400 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 6888 0 6944 400 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 30968 0 31024 400 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 9128 0 9184 400 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 10808 0 10864 400 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 12488 0 12544 400 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 15288 0 15344 400 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 16968 0 17024 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 17808 0 17864 400 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 18648 0 18704 400 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 20328 0 20384 400 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 22008 0 22064 400 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 23688 0 23744 400 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 24528 0 24584 400 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 25368 0 25424 400 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 26208 0 26264 400 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 27048 0 27104 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 28728 0 28784 400 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 30408 0 30464 400 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 31248 0 31304 400 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 32088 0 32144 400 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 10248 0 10304 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 11088 0 11144 400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 11928 0 11984 400 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 12768 0 12824 400 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 13608 0 13664 400 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 5208 0 5264 400 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 14728 0 14784 400 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 16408 0 16464 400 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 18088 0 18144 400 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 19768 0 19824 400 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 21448 0 21504 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 6328 0 6384 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 23128 0 23184 400 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 24808 0 24864 400 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 26488 0 26544 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 27328 0 27384 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 29848 0 29904 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 7448 0 7504 400 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 31528 0 31584 400 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 8568 0 8624 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 9688 0 9744 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 11368 0 11424 400 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 13048 0 13104 400 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 13888 0 13944 400 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 5488 0 5544 400 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 4088 0 4144 400 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3433480
string GDS_FILE /home/rs2xd/gf180_shuttle/gf180-demo/openlane/user_proj_example/runs/22_11_30_09_32/results/signoff/user_proj_example.magic.gds
string GDS_START 200846
<< end >>

