magic
tech gf180mcuC
magscale 1 5
timestamp 1670096991
<< metal2 >>
rect 5796 299760 5908 300480
rect 16884 299796 16996 300480
rect 16870 299760 16996 299796
rect 27734 299782 27930 299810
rect 27972 299796 28084 300480
rect 15526 297906 15554 297911
rect 2086 295722 2114 295727
rect 2086 257474 2114 295694
rect 10038 289842 10066 289847
rect 5446 288610 5474 288615
rect 2086 257441 2114 257446
rect 3766 274386 3794 274391
rect 2198 255906 2226 255911
rect 2142 255122 2170 255127
rect 2086 245714 2114 245719
rect 2086 182042 2114 245686
rect 2142 210490 2170 255094
rect 2198 231826 2226 255878
rect 2198 231793 2226 231798
rect 2142 210457 2170 210462
rect 2198 224602 2226 224607
rect 2086 182009 2114 182014
rect 2086 139258 2114 139263
rect 2086 32354 2114 139230
rect 2198 139034 2226 224574
rect 2198 139001 2226 139006
rect 2086 32321 2114 32326
rect 2142 125034 2170 125039
rect 2142 31906 2170 125006
rect 2310 61026 2338 61031
rect 2310 54194 2338 60998
rect 2310 54161 2338 54166
rect 2142 31873 2170 31878
rect 2198 53914 2226 53919
rect 2198 15554 2226 53886
rect 2310 39690 2338 39695
rect 2310 36106 2338 39662
rect 3766 39522 3794 274358
rect 5446 259154 5474 288582
rect 5446 259121 5474 259126
rect 7966 267162 7994 267167
rect 6286 256410 6314 256415
rect 5446 255514 5474 255519
rect 3766 39489 3794 39494
rect 3822 189042 3850 189047
rect 2310 36073 2338 36078
rect 2926 32354 2954 32359
rect 2926 24346 2954 32326
rect 3262 31906 3290 31911
rect 3262 29834 3290 31878
rect 3262 29801 3290 29806
rect 2926 24313 2954 24318
rect 3766 24346 3794 24351
rect 3766 21434 3794 24318
rect 3766 21401 3794 21406
rect 2198 15521 2226 15526
rect 3822 14322 3850 189014
rect 5446 167818 5474 255486
rect 5446 167785 5474 167790
rect 5894 221802 5922 221807
rect 5502 155442 5530 155447
rect 5446 146370 5474 146375
rect 4606 36106 4634 36111
rect 4606 33138 4634 36078
rect 4606 33105 4634 33110
rect 5054 33138 5082 33143
rect 5054 30674 5082 33110
rect 5054 30641 5082 30646
rect 5446 14378 5474 146342
rect 5502 103810 5530 155414
rect 5502 103777 5530 103782
rect 5446 14345 5474 14350
rect 3822 14289 3850 14294
rect 5894 210 5922 221774
rect 6286 203322 6314 256382
rect 7182 256298 7210 256303
rect 7126 252882 7154 252887
rect 7126 237762 7154 252854
rect 7126 237729 7154 237734
rect 6286 203289 6314 203294
rect 7126 196602 7154 196607
rect 6846 30674 6874 30679
rect 6846 30058 6874 30646
rect 6846 30025 6874 30030
rect 6286 29834 6314 29839
rect 6286 26922 6314 29806
rect 6286 26889 6314 26894
rect 6958 21434 6986 21439
rect 6958 18074 6986 21406
rect 6958 18041 6986 18046
rect 7126 17682 7154 196574
rect 7182 160482 7210 256270
rect 7182 160449 7210 160454
rect 7966 31122 7994 267134
rect 8918 256466 8946 256471
rect 8862 246162 8890 246167
rect 8806 245322 8834 245327
rect 7966 31089 7994 31094
rect 8022 139034 8050 139039
rect 7966 30058 7994 30063
rect 7966 27762 7994 30030
rect 7966 27729 7994 27734
rect 7126 17649 7154 17654
rect 8022 14266 8050 139006
rect 8022 14233 8050 14238
rect 8806 14210 8834 245294
rect 8862 117642 8890 246134
rect 8918 245714 8946 256438
rect 8918 245681 8946 245686
rect 8862 117609 8890 117614
rect 8862 27762 8890 27767
rect 8862 20986 8890 27734
rect 9254 26866 9282 26871
rect 9254 25186 9282 26838
rect 9254 25153 9282 25158
rect 10038 22722 10066 289814
rect 14630 261674 14658 261679
rect 10878 260050 10906 260055
rect 10038 22689 10066 22694
rect 10486 74802 10514 74807
rect 8862 20953 8890 20958
rect 10486 14490 10514 74774
rect 10878 47922 10906 260022
rect 12558 259994 12586 259999
rect 12502 255234 12530 255239
rect 12502 147434 12530 255206
rect 12502 147401 12530 147406
rect 10878 47889 10906 47894
rect 12166 89250 12194 89255
rect 12166 31962 12194 89222
rect 12558 56378 12586 259966
rect 14294 258370 14322 258375
rect 13342 258314 13370 258319
rect 13342 139034 13370 258286
rect 14182 255682 14210 255687
rect 13342 139001 13370 139006
rect 13398 255178 13426 255183
rect 12558 56345 12586 56350
rect 12166 31929 12194 31934
rect 12222 54194 12250 54199
rect 10934 25186 10962 25191
rect 10934 23954 10962 25158
rect 10934 23921 10962 23926
rect 10934 20986 10962 20991
rect 10934 19754 10962 20958
rect 10934 19721 10962 19726
rect 12166 19754 12194 19759
rect 12166 18522 12194 19726
rect 12166 18489 12194 18494
rect 10486 14457 10514 14462
rect 8806 14177 8834 14182
rect 12222 14154 12250 54166
rect 13006 23954 13034 23959
rect 13006 21042 13034 23926
rect 13006 21009 13034 21014
rect 13398 15946 13426 255150
rect 14126 251202 14154 251207
rect 14126 188762 14154 251174
rect 14126 188729 14154 188734
rect 14182 163898 14210 255654
rect 14182 163865 14210 163870
rect 14238 252042 14266 252047
rect 13454 97650 13482 97655
rect 13454 96642 13482 97622
rect 13454 96609 13482 96614
rect 14238 81242 14266 252014
rect 14238 81209 14266 81214
rect 14238 72786 14266 72791
rect 13902 21042 13930 21047
rect 13902 19306 13930 21014
rect 13902 19273 13930 19278
rect 14238 16002 14266 72758
rect 14294 64442 14322 258342
rect 14462 255850 14490 255855
rect 14350 255794 14378 255799
rect 14350 180698 14378 255766
rect 14462 230426 14490 255822
rect 14462 230393 14490 230398
rect 14350 180665 14378 180670
rect 14294 64409 14322 64414
rect 14350 106050 14378 106055
rect 14238 15974 14322 16002
rect 13398 15913 13426 15918
rect 12222 14121 12250 14126
rect 14294 13986 14322 15974
rect 14350 14826 14378 106022
rect 14350 14793 14378 14798
rect 14294 13953 14322 13958
rect 7574 13874 7602 13879
rect 6566 240 6650 266
rect 7574 240 7602 13846
rect 14630 13370 14658 261646
rect 14686 257082 14714 257087
rect 14686 252042 14714 257054
rect 15526 255178 15554 297878
rect 16366 297794 16394 297799
rect 16366 255682 16394 297766
rect 16870 294014 16898 299760
rect 16814 293986 16898 294014
rect 16814 259210 16842 293986
rect 23646 275114 23674 275119
rect 21014 272594 21042 272599
rect 19726 271418 19754 271423
rect 18494 268002 18522 268007
rect 18494 266322 18522 267974
rect 19726 268002 19754 271390
rect 21014 271418 21042 272566
rect 23646 272594 23674 275086
rect 23646 272561 23674 272566
rect 21014 271385 21042 271390
rect 19726 267969 19754 267974
rect 18438 266294 18522 266322
rect 17206 265874 17234 265879
rect 17206 261674 17234 265846
rect 18438 265874 18466 266294
rect 18438 265841 18466 265846
rect 17206 261641 17234 261646
rect 16814 259177 16842 259182
rect 16366 255649 16394 255654
rect 23086 256578 23114 256583
rect 15526 255145 15554 255150
rect 23086 254884 23114 256550
rect 27734 255850 27762 299782
rect 27902 299754 27930 299782
rect 27958 299760 28084 299796
rect 39060 299760 39172 300480
rect 50148 299796 50260 300480
rect 50134 299760 50260 299796
rect 60494 299782 61194 299810
rect 61236 299796 61348 300480
rect 27958 299754 27986 299760
rect 27902 299726 27986 299754
rect 32326 297850 32354 297855
rect 27734 255817 27762 255822
rect 31486 256746 31514 256751
rect 31486 254884 31514 256718
rect 32326 256746 32354 297822
rect 50134 297850 50162 299760
rect 50134 297817 50162 297822
rect 57134 281834 57162 281839
rect 52486 279314 52514 279319
rect 52486 275114 52514 279286
rect 57134 279314 57162 281806
rect 57134 279281 57162 279286
rect 52486 275081 52514 275086
rect 32326 256713 32354 256718
rect 39550 256354 39578 256359
rect 39550 254884 39578 256326
rect 60494 255794 60522 299782
rect 61166 299754 61194 299782
rect 61222 299760 61348 299796
rect 72324 299760 72436 300480
rect 83174 299782 83370 299810
rect 83412 299796 83524 300480
rect 61222 299754 61250 299760
rect 61166 299726 61250 299754
rect 80206 288554 80234 288559
rect 80206 281834 80234 288526
rect 83174 288554 83202 299782
rect 83342 299754 83370 299782
rect 83398 299760 83524 299796
rect 94500 299796 94612 300480
rect 94500 299760 94626 299796
rect 105588 299760 105700 300480
rect 116676 299796 116788 300480
rect 127764 299796 127876 300480
rect 116662 299760 116788 299796
rect 127750 299760 127876 299796
rect 138852 299760 138964 300480
rect 149534 299782 149898 299810
rect 149940 299796 150052 300480
rect 83398 299754 83426 299760
rect 83342 299726 83426 299754
rect 94598 297850 94626 299760
rect 116662 297906 116690 299760
rect 116662 297873 116690 297878
rect 94598 297817 94626 297822
rect 127750 294014 127778 299760
rect 83174 288521 83202 288526
rect 127694 293986 127778 294014
rect 80206 281801 80234 281806
rect 105854 259210 105882 259215
rect 97678 257530 97706 257535
rect 60494 255761 60522 255766
rect 61670 256354 61698 256359
rect 61670 255794 61698 256326
rect 61670 255761 61698 255766
rect 64414 256354 64442 256359
rect 64414 254884 64442 256326
rect 89278 255458 89306 255463
rect 89278 254884 89306 255430
rect 97678 254884 97706 257502
rect 105854 254898 105882 259182
rect 127694 255850 127722 293986
rect 149534 258370 149562 299782
rect 149870 299754 149898 299782
rect 149926 299760 150052 299796
rect 160454 299782 160986 299810
rect 161028 299796 161140 300480
rect 149926 299754 149954 299760
rect 149870 299726 149954 299754
rect 160454 260050 160482 299782
rect 160958 299754 160986 299782
rect 161014 299760 161140 299796
rect 172116 299760 172228 300480
rect 183204 299796 183316 300480
rect 194292 299796 194404 300480
rect 183204 299760 183330 299796
rect 194292 299760 194418 299796
rect 205380 299760 205492 300480
rect 216468 299796 216580 300480
rect 216468 299760 216594 299796
rect 161014 299754 161042 299760
rect 160958 299726 161042 299754
rect 183302 294434 183330 299760
rect 194390 295946 194418 299760
rect 216566 297906 216594 299760
rect 216566 297873 216594 297878
rect 226814 299782 227514 299810
rect 227556 299796 227668 300480
rect 221326 297850 221354 297855
rect 194390 295913 194418 295918
rect 196126 295946 196154 295951
rect 183302 294401 183330 294406
rect 188566 294434 188594 294439
rect 188566 283906 188594 294406
rect 196126 291354 196154 295918
rect 196126 291321 196154 291326
rect 199486 291354 199514 291359
rect 199486 287714 199514 291326
rect 199486 287681 199514 287686
rect 201166 287714 201194 287719
rect 188566 283873 188594 283878
rect 190246 283906 190274 283911
rect 190246 268394 190274 283878
rect 201166 280602 201194 287686
rect 201166 280569 201194 280574
rect 204134 280602 204162 280607
rect 204134 278474 204162 280574
rect 204134 278441 204162 278446
rect 206206 278474 206234 278479
rect 206206 275954 206234 278446
rect 206206 275921 206234 275926
rect 219534 275954 219562 275959
rect 219534 271754 219562 275926
rect 219534 271721 219562 271726
rect 190246 268361 190274 268366
rect 196966 268394 196994 268399
rect 160454 260017 160482 260022
rect 180614 259154 180642 259159
rect 180614 258734 180642 259126
rect 180614 258706 180698 258734
rect 149534 258337 149562 258342
rect 155806 256522 155834 256527
rect 127694 255817 127722 255822
rect 130550 255906 130578 255911
rect 122150 255514 122178 255519
rect 122150 254898 122178 255486
rect 130550 254898 130578 255878
rect 147406 255514 147434 255519
rect 105854 254870 106036 254898
rect 122150 254870 122500 254898
rect 130550 254870 130900 254898
rect 147406 254884 147434 255486
rect 155806 254884 155834 256494
rect 163870 256466 163898 256471
rect 163870 254884 163898 256438
rect 172270 255570 172298 255575
rect 172270 254884 172298 255542
rect 180670 254884 180698 258706
rect 196966 258482 196994 268366
rect 196966 258449 196994 258454
rect 188734 258370 188762 258375
rect 188734 254884 188762 258342
rect 221326 257138 221354 297822
rect 226366 271754 226394 271759
rect 226366 265034 226394 271726
rect 226366 265001 226394 265006
rect 226814 257530 226842 299782
rect 227486 299754 227514 299782
rect 227542 299760 227668 299796
rect 238644 299760 238756 300480
rect 249494 299782 249690 299810
rect 249732 299796 249844 300480
rect 227542 299754 227570 299760
rect 227486 299726 227570 299754
rect 233086 265034 233114 265039
rect 233086 262514 233114 265006
rect 233086 262481 233114 262486
rect 236614 262514 236642 262519
rect 236614 260386 236642 262486
rect 236614 260353 236642 260358
rect 238966 260386 238994 260391
rect 231798 258482 231826 258487
rect 226814 257497 226842 257502
rect 230398 258426 230426 258431
rect 221326 257105 221354 257110
rect 221774 257138 221802 257143
rect 197134 256466 197162 256471
rect 197134 254884 197162 256438
rect 213374 256410 213402 256415
rect 213374 254898 213402 256382
rect 221774 254898 221802 257110
rect 213374 254870 213556 254898
rect 221774 254870 221956 254898
rect 230398 254884 230426 258398
rect 231798 257530 231826 258454
rect 231798 257497 231826 257502
rect 238966 256634 238994 260358
rect 238966 256601 238994 256606
rect 238070 256298 238098 256303
rect 238070 254898 238098 256270
rect 249494 255906 249522 299782
rect 249662 299754 249690 299782
rect 249718 299760 249844 299796
rect 260414 299782 260778 299810
rect 260820 299796 260932 300480
rect 249718 299754 249746 299760
rect 249662 299726 249746 299754
rect 255486 297906 255514 297911
rect 255150 257530 255178 257535
rect 249494 255873 249522 255878
rect 255038 257082 255066 257087
rect 238070 254870 238420 254898
rect 14686 252009 14714 252014
rect 14742 253666 14770 253671
rect 14742 251202 14770 253638
rect 14742 251169 14770 251174
rect 255038 224266 255066 257054
rect 255038 224233 255066 224238
rect 14686 82362 14714 82372
rect 14686 14434 14714 82334
rect 255094 42770 255122 42775
rect 254982 39578 255010 39583
rect 14686 14401 14714 14406
rect 14742 19306 14770 19311
rect 14742 13426 14770 19278
rect 14910 18466 14938 18471
rect 14798 18074 14826 18079
rect 14798 14938 14826 18046
rect 14798 14905 14826 14910
rect 14910 14882 14938 18438
rect 14966 15946 14994 15951
rect 14966 15372 14994 15918
rect 14910 14849 14938 14854
rect 15246 15106 15274 15111
rect 15246 14098 15274 15078
rect 23030 14266 23058 15148
rect 23030 14233 23058 14238
rect 56294 14210 56322 15148
rect 64358 14490 64386 15148
rect 64358 14457 64386 14462
rect 72758 14434 72786 15148
rect 72758 14401 72786 14406
rect 56294 14177 56322 14182
rect 81214 14210 81242 15148
rect 81214 14177 81242 14182
rect 15246 14065 15274 14070
rect 97622 14098 97650 15148
rect 106022 14154 106050 15148
rect 106022 14121 106050 14126
rect 97622 14065 97650 14070
rect 130942 14098 130970 15148
rect 130942 14065 130970 14070
rect 14742 13393 14770 13398
rect 14630 13337 14658 13342
rect 139006 13314 139034 15148
rect 147406 14154 147434 15148
rect 163814 14378 163842 15148
rect 163814 14345 163842 14350
rect 166110 14714 166138 14719
rect 147406 14121 147434 14126
rect 166110 14098 166138 14686
rect 166110 14065 166138 14070
rect 172214 13370 172242 15148
rect 180670 14098 180698 15148
rect 197134 14378 197162 15148
rect 197134 14345 197162 14350
rect 180670 14065 180698 14070
rect 221998 14042 222026 15148
rect 246806 14322 246834 15148
rect 254982 14882 255010 39550
rect 254982 14849 255010 14854
rect 255038 25914 255066 25919
rect 246806 14289 246834 14294
rect 221998 14009 222026 14014
rect 255038 13986 255066 25886
rect 255094 14938 255122 42742
rect 255094 14905 255122 14910
rect 255038 13953 255066 13958
rect 172214 13337 172242 13342
rect 139006 13281 139034 13286
rect 255150 13314 255178 257502
rect 255374 255906 255402 255911
rect 255374 14042 255402 255878
rect 255430 255850 255458 255855
rect 255430 23114 255458 255822
rect 255486 205562 255514 297878
rect 258286 283122 258314 283127
rect 258286 258370 258314 283094
rect 260414 259994 260442 299782
rect 260750 299754 260778 299782
rect 260806 299760 260932 299796
rect 271908 299760 272020 300480
rect 282996 299796 283108 300480
rect 294084 299796 294196 300480
rect 282982 299760 283108 299796
rect 294070 299760 294196 299796
rect 260806 299754 260834 299760
rect 260750 299726 260834 299754
rect 260414 259961 260442 259966
rect 275086 297850 275114 297855
rect 258286 258337 258314 258342
rect 257054 257474 257082 257479
rect 256606 224266 256634 224271
rect 256606 219674 256634 224238
rect 256606 219641 256634 219646
rect 255486 205529 255514 205534
rect 255430 23081 255458 23086
rect 255766 139034 255794 139039
rect 255374 14009 255402 14014
rect 255766 13426 255794 139006
rect 257054 122570 257082 257446
rect 258286 256522 258314 256527
rect 257110 255122 257138 255127
rect 257110 238490 257138 255094
rect 257110 238457 257138 238462
rect 257446 246890 257474 246895
rect 257054 122537 257082 122542
rect 257110 130970 257138 130975
rect 256662 114170 256690 114175
rect 256662 113442 256690 114142
rect 256662 113409 256690 113414
rect 256214 47978 256242 47983
rect 256214 42770 256242 47950
rect 256214 42737 256242 42742
rect 256606 29834 256634 29839
rect 256606 25914 256634 29806
rect 256606 25881 256634 25886
rect 257110 13874 257138 130942
rect 257110 13841 257138 13846
rect 255766 13393 255794 13398
rect 255150 13281 255178 13286
rect 257446 3402 257474 246862
rect 258286 164234 258314 256494
rect 262486 255570 262514 255575
rect 260862 255402 260890 255407
rect 260806 249522 260834 249527
rect 258286 164201 258314 164206
rect 259126 230202 259154 230207
rect 257894 163898 257922 163903
rect 257894 10962 257922 163870
rect 258286 147434 258314 147439
rect 258286 103362 258314 147406
rect 258286 103329 258314 103334
rect 258286 89306 258314 89311
rect 258286 42882 258314 89278
rect 258286 42849 258314 42854
rect 259126 22722 259154 230174
rect 260806 56322 260834 249494
rect 260862 248234 260890 255374
rect 260862 248201 260890 248206
rect 262486 183162 262514 255542
rect 267526 255514 267554 255519
rect 266686 255458 266714 255463
rect 265846 248234 265874 248239
rect 265846 245714 265874 248206
rect 265846 245681 265874 245686
rect 262486 183129 262514 183134
rect 261646 97482 261674 97487
rect 261646 83202 261674 97454
rect 261646 83169 261674 83174
rect 260806 56289 260834 56294
rect 261646 69762 261674 69767
rect 260806 34874 260834 34879
rect 260806 29834 260834 34846
rect 260806 29801 260834 29806
rect 259126 22689 259154 22694
rect 261646 14154 261674 69734
rect 266686 63042 266714 255430
rect 267526 122682 267554 255486
rect 270606 245714 270634 245719
rect 270606 243194 270634 245686
rect 270606 243161 270634 243166
rect 274246 219674 274274 219679
rect 274246 212954 274274 219646
rect 274246 212921 274274 212926
rect 267526 122649 267554 122654
rect 268366 209202 268394 209207
rect 266686 63009 266714 63014
rect 265846 39522 265874 39527
rect 265846 34874 265874 39494
rect 265846 34841 265874 34846
rect 268366 14378 268394 209174
rect 275086 188202 275114 297822
rect 282982 297850 283010 299760
rect 282982 297817 283010 297822
rect 294070 297794 294098 299760
rect 294070 297761 294098 297766
rect 297766 269906 297794 269911
rect 282646 262962 282674 262967
rect 282646 258426 282674 262934
rect 282646 258393 282674 258398
rect 297766 258314 297794 269878
rect 297766 258281 297794 258286
rect 275086 188169 275114 188174
rect 279286 256578 279314 256583
rect 279286 129402 279314 256550
rect 280126 256466 280154 256471
rect 279342 243194 279370 243199
rect 279342 239834 279370 243166
rect 279342 239801 279370 239806
rect 279286 129369 279314 129374
rect 280126 109242 280154 256438
rect 282646 256354 282674 256359
rect 280182 212954 280210 212959
rect 280182 209594 280210 212926
rect 280182 209561 280210 209566
rect 280126 109209 280154 109214
rect 280966 203322 280994 203327
rect 276766 105882 276794 105892
rect 275926 77714 275954 77719
rect 273742 51282 273770 51287
rect 271726 48706 271754 48711
rect 270046 42434 270074 42439
rect 270046 39522 270074 42406
rect 271726 42434 271754 48678
rect 273742 48706 273770 51254
rect 275926 51282 275954 77686
rect 275926 51249 275954 51254
rect 273742 48673 273770 48678
rect 271726 42401 271754 42406
rect 270046 39489 270074 39494
rect 268366 14345 268394 14350
rect 261646 14121 261674 14126
rect 257894 10929 257922 10934
rect 276766 9282 276794 105854
rect 280574 81074 280602 81079
rect 280574 77714 280602 81046
rect 280574 77681 280602 77686
rect 280966 72282 280994 203294
rect 282646 149562 282674 256326
rect 297766 255794 297794 255799
rect 297766 223370 297794 255766
rect 297822 255178 297850 255183
rect 297822 243362 297850 255150
rect 297822 243329 297850 243334
rect 297822 239834 297850 239839
rect 297822 230034 297850 239806
rect 297822 230001 297850 230006
rect 297766 223337 297794 223342
rect 284326 209594 284354 209599
rect 284326 200746 284354 209566
rect 284326 200713 284354 200718
rect 286846 200746 286874 200751
rect 286846 194474 286874 200718
rect 286846 194441 286874 194446
rect 290206 194474 290234 194479
rect 290206 192402 290234 194446
rect 290206 192369 290234 192374
rect 292110 192402 292138 192407
rect 292110 189882 292138 192374
rect 292110 189849 292138 189854
rect 282646 149529 282674 149534
rect 288526 169722 288554 169727
rect 280966 72249 280994 72254
rect 288526 14098 288554 169694
rect 297374 164234 297402 164239
rect 297374 163394 297402 164206
rect 297374 163361 297402 163366
rect 297766 143290 297794 143295
rect 297766 113442 297794 143262
rect 297766 113409 297794 113414
rect 290206 89922 290234 89927
rect 290206 81074 290234 89894
rect 290206 81041 290234 81046
rect 297766 49994 297794 49999
rect 297766 14714 297794 49966
rect 297878 30002 297906 30007
rect 297878 14826 297906 29974
rect 297878 14793 297906 14798
rect 297766 14681 297794 14686
rect 288526 14065 288554 14070
rect 276766 9249 276794 9254
rect 257446 3369 257474 3374
rect 6566 238 6748 240
rect 6566 210 6594 238
rect 5894 182 6594 210
rect 6622 196 6748 238
rect 7574 196 7700 240
rect 6636 -480 6748 196
rect 7588 -480 7700 196
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
rect 293188 -480 293300 240
<< via2 >>
rect 15526 297878 15554 297906
rect 2086 295694 2114 295722
rect 10038 289814 10066 289842
rect 5446 288582 5474 288610
rect 2086 257446 2114 257474
rect 3766 274358 3794 274386
rect 2198 255878 2226 255906
rect 2142 255094 2170 255122
rect 2086 245686 2114 245714
rect 2198 231798 2226 231826
rect 2142 210462 2170 210490
rect 2198 224574 2226 224602
rect 2086 182014 2114 182042
rect 2086 139230 2114 139258
rect 2198 139006 2226 139034
rect 2086 32326 2114 32354
rect 2142 125006 2170 125034
rect 2310 60998 2338 61026
rect 2310 54166 2338 54194
rect 2142 31878 2170 31906
rect 2198 53886 2226 53914
rect 2310 39662 2338 39690
rect 5446 259126 5474 259154
rect 7966 267134 7994 267162
rect 6286 256382 6314 256410
rect 5446 255486 5474 255514
rect 3766 39494 3794 39522
rect 3822 189014 3850 189042
rect 2310 36078 2338 36106
rect 2926 32326 2954 32354
rect 3262 31878 3290 31906
rect 3262 29806 3290 29834
rect 2926 24318 2954 24346
rect 3766 24318 3794 24346
rect 3766 21406 3794 21434
rect 2198 15526 2226 15554
rect 5446 167790 5474 167818
rect 5894 221774 5922 221802
rect 5502 155414 5530 155442
rect 5446 146342 5474 146370
rect 4606 36078 4634 36106
rect 4606 33110 4634 33138
rect 5054 33110 5082 33138
rect 5054 30646 5082 30674
rect 5502 103782 5530 103810
rect 5446 14350 5474 14378
rect 3822 14294 3850 14322
rect 7182 256270 7210 256298
rect 7126 252854 7154 252882
rect 7126 237734 7154 237762
rect 6286 203294 6314 203322
rect 7126 196574 7154 196602
rect 6846 30646 6874 30674
rect 6846 30030 6874 30058
rect 6286 29806 6314 29834
rect 6286 26894 6314 26922
rect 6958 21406 6986 21434
rect 6958 18046 6986 18074
rect 7182 160454 7210 160482
rect 8918 256438 8946 256466
rect 8862 246134 8890 246162
rect 8806 245294 8834 245322
rect 7966 31094 7994 31122
rect 8022 139006 8050 139034
rect 7966 30030 7994 30058
rect 7966 27734 7994 27762
rect 7126 17654 7154 17682
rect 8022 14238 8050 14266
rect 8918 245686 8946 245714
rect 8862 117614 8890 117642
rect 8862 27734 8890 27762
rect 9254 26838 9282 26866
rect 9254 25158 9282 25186
rect 14630 261646 14658 261674
rect 10878 260022 10906 260050
rect 10038 22694 10066 22722
rect 10486 74774 10514 74802
rect 8862 20958 8890 20986
rect 12558 259966 12586 259994
rect 12502 255206 12530 255234
rect 12502 147406 12530 147434
rect 10878 47894 10906 47922
rect 12166 89222 12194 89250
rect 14294 258342 14322 258370
rect 13342 258286 13370 258314
rect 14182 255654 14210 255682
rect 13342 139006 13370 139034
rect 13398 255150 13426 255178
rect 12558 56350 12586 56378
rect 12166 31934 12194 31962
rect 12222 54166 12250 54194
rect 10934 25158 10962 25186
rect 10934 23926 10962 23954
rect 10934 20958 10962 20986
rect 10934 19726 10962 19754
rect 12166 19726 12194 19754
rect 12166 18494 12194 18522
rect 10486 14462 10514 14490
rect 8806 14182 8834 14210
rect 13006 23926 13034 23954
rect 13006 21014 13034 21042
rect 14126 251174 14154 251202
rect 14126 188734 14154 188762
rect 14182 163870 14210 163898
rect 14238 252014 14266 252042
rect 13454 97622 13482 97650
rect 13454 96614 13482 96642
rect 14238 81214 14266 81242
rect 14238 72758 14266 72786
rect 13902 21014 13930 21042
rect 13902 19278 13930 19306
rect 14462 255822 14490 255850
rect 14350 255766 14378 255794
rect 14462 230398 14490 230426
rect 14350 180670 14378 180698
rect 14294 64414 14322 64442
rect 14350 106022 14378 106050
rect 13398 15918 13426 15946
rect 12222 14126 12250 14154
rect 14350 14798 14378 14826
rect 14294 13958 14322 13986
rect 7574 13846 7602 13874
rect 14686 257054 14714 257082
rect 16366 297766 16394 297794
rect 23646 275086 23674 275114
rect 21014 272566 21042 272594
rect 19726 271390 19754 271418
rect 18494 267974 18522 268002
rect 23646 272566 23674 272594
rect 21014 271390 21042 271418
rect 19726 267974 19754 268002
rect 17206 265846 17234 265874
rect 18438 265846 18466 265874
rect 17206 261646 17234 261674
rect 16814 259182 16842 259210
rect 16366 255654 16394 255682
rect 23086 256550 23114 256578
rect 15526 255150 15554 255178
rect 32326 297822 32354 297850
rect 27734 255822 27762 255850
rect 31486 256718 31514 256746
rect 50134 297822 50162 297850
rect 57134 281806 57162 281834
rect 52486 279286 52514 279314
rect 57134 279286 57162 279314
rect 52486 275086 52514 275114
rect 32326 256718 32354 256746
rect 39550 256326 39578 256354
rect 80206 288526 80234 288554
rect 116662 297878 116690 297906
rect 94598 297822 94626 297850
rect 83174 288526 83202 288554
rect 80206 281806 80234 281834
rect 105854 259182 105882 259210
rect 97678 257502 97706 257530
rect 60494 255766 60522 255794
rect 61670 256326 61698 256354
rect 61670 255766 61698 255794
rect 64414 256326 64442 256354
rect 89278 255430 89306 255458
rect 216566 297878 216594 297906
rect 221326 297822 221354 297850
rect 194390 295918 194418 295946
rect 196126 295918 196154 295946
rect 183302 294406 183330 294434
rect 188566 294406 188594 294434
rect 196126 291326 196154 291354
rect 199486 291326 199514 291354
rect 199486 287686 199514 287714
rect 201166 287686 201194 287714
rect 188566 283878 188594 283906
rect 190246 283878 190274 283906
rect 201166 280574 201194 280602
rect 204134 280574 204162 280602
rect 204134 278446 204162 278474
rect 206206 278446 206234 278474
rect 206206 275926 206234 275954
rect 219534 275926 219562 275954
rect 219534 271726 219562 271754
rect 190246 268366 190274 268394
rect 196966 268366 196994 268394
rect 160454 260022 160482 260050
rect 180614 259126 180642 259154
rect 149534 258342 149562 258370
rect 155806 256494 155834 256522
rect 127694 255822 127722 255850
rect 130550 255878 130578 255906
rect 122150 255486 122178 255514
rect 147406 255486 147434 255514
rect 163870 256438 163898 256466
rect 172270 255542 172298 255570
rect 196966 258454 196994 258482
rect 188734 258342 188762 258370
rect 226366 271726 226394 271754
rect 226366 265006 226394 265034
rect 233086 265006 233114 265034
rect 233086 262486 233114 262514
rect 236614 262486 236642 262514
rect 236614 260358 236642 260386
rect 238966 260358 238994 260386
rect 231798 258454 231826 258482
rect 226814 257502 226842 257530
rect 230398 258398 230426 258426
rect 221326 257110 221354 257138
rect 221774 257110 221802 257138
rect 197134 256438 197162 256466
rect 213374 256382 213402 256410
rect 231798 257502 231826 257530
rect 238966 256606 238994 256634
rect 238070 256270 238098 256298
rect 255486 297878 255514 297906
rect 255150 257502 255178 257530
rect 249494 255878 249522 255906
rect 255038 257054 255066 257082
rect 14686 252014 14714 252042
rect 14742 253638 14770 253666
rect 14742 251174 14770 251202
rect 255038 224238 255066 224266
rect 14686 82334 14714 82362
rect 255094 42742 255122 42770
rect 254982 39550 255010 39578
rect 14686 14406 14714 14434
rect 14742 19278 14770 19306
rect 14910 18438 14938 18466
rect 14798 18046 14826 18074
rect 14798 14910 14826 14938
rect 14966 15918 14994 15946
rect 14910 14854 14938 14882
rect 15246 15078 15274 15106
rect 23030 14238 23058 14266
rect 64358 14462 64386 14490
rect 72758 14406 72786 14434
rect 56294 14182 56322 14210
rect 81214 14182 81242 14210
rect 15246 14070 15274 14098
rect 106022 14126 106050 14154
rect 97622 14070 97650 14098
rect 130942 14070 130970 14098
rect 14742 13398 14770 13426
rect 14630 13342 14658 13370
rect 163814 14350 163842 14378
rect 166110 14686 166138 14714
rect 147406 14126 147434 14154
rect 166110 14070 166138 14098
rect 197134 14350 197162 14378
rect 180670 14070 180698 14098
rect 254982 14854 255010 14882
rect 255038 25886 255066 25914
rect 246806 14294 246834 14322
rect 221998 14014 222026 14042
rect 255094 14910 255122 14938
rect 255038 13958 255066 13986
rect 172214 13342 172242 13370
rect 139006 13286 139034 13314
rect 255374 255878 255402 255906
rect 255430 255822 255458 255850
rect 258286 283094 258314 283122
rect 260414 259966 260442 259994
rect 275086 297822 275114 297850
rect 258286 258342 258314 258370
rect 257054 257446 257082 257474
rect 256606 224238 256634 224266
rect 256606 219646 256634 219674
rect 255486 205534 255514 205562
rect 255430 23086 255458 23114
rect 255766 139006 255794 139034
rect 255374 14014 255402 14042
rect 258286 256494 258314 256522
rect 257110 255094 257138 255122
rect 257110 238462 257138 238490
rect 257446 246862 257474 246890
rect 257054 122542 257082 122570
rect 257110 130942 257138 130970
rect 256662 114142 256690 114170
rect 256662 113414 256690 113442
rect 256214 47950 256242 47978
rect 256214 42742 256242 42770
rect 256606 29806 256634 29834
rect 256606 25886 256634 25914
rect 257110 13846 257138 13874
rect 255766 13398 255794 13426
rect 255150 13286 255178 13314
rect 262486 255542 262514 255570
rect 260862 255374 260890 255402
rect 260806 249494 260834 249522
rect 258286 164206 258314 164234
rect 259126 230174 259154 230202
rect 257894 163870 257922 163898
rect 258286 147406 258314 147434
rect 258286 103334 258314 103362
rect 258286 89278 258314 89306
rect 258286 42854 258314 42882
rect 260862 248206 260890 248234
rect 267526 255486 267554 255514
rect 266686 255430 266714 255458
rect 265846 248206 265874 248234
rect 265846 245686 265874 245714
rect 262486 183134 262514 183162
rect 261646 97454 261674 97482
rect 261646 83174 261674 83202
rect 260806 56294 260834 56322
rect 261646 69734 261674 69762
rect 260806 34846 260834 34874
rect 260806 29806 260834 29834
rect 259126 22694 259154 22722
rect 270606 245686 270634 245714
rect 270606 243166 270634 243194
rect 274246 219646 274274 219674
rect 274246 212926 274274 212954
rect 267526 122654 267554 122682
rect 268366 209174 268394 209202
rect 266686 63014 266714 63042
rect 265846 39494 265874 39522
rect 265846 34846 265874 34874
rect 282982 297822 283010 297850
rect 294070 297766 294098 297794
rect 297766 269878 297794 269906
rect 282646 262934 282674 262962
rect 282646 258398 282674 258426
rect 297766 258286 297794 258314
rect 275086 188174 275114 188202
rect 279286 256550 279314 256578
rect 280126 256438 280154 256466
rect 279342 243166 279370 243194
rect 279342 239806 279370 239834
rect 279286 129374 279314 129402
rect 282646 256326 282674 256354
rect 280182 212926 280210 212954
rect 280182 209566 280210 209594
rect 280126 109214 280154 109242
rect 280966 203294 280994 203322
rect 276766 105854 276794 105882
rect 275926 77686 275954 77714
rect 273742 51254 273770 51282
rect 271726 48678 271754 48706
rect 270046 42406 270074 42434
rect 275926 51254 275954 51282
rect 273742 48678 273770 48706
rect 271726 42406 271754 42434
rect 270046 39494 270074 39522
rect 268366 14350 268394 14378
rect 261646 14126 261674 14154
rect 257894 10934 257922 10962
rect 280574 81046 280602 81074
rect 280574 77686 280602 77714
rect 297766 255766 297794 255794
rect 297822 255150 297850 255178
rect 297822 243334 297850 243362
rect 297822 239806 297850 239834
rect 297822 230006 297850 230034
rect 297766 223342 297794 223370
rect 284326 209566 284354 209594
rect 284326 200718 284354 200746
rect 286846 200718 286874 200746
rect 286846 194446 286874 194474
rect 290206 194446 290234 194474
rect 290206 192374 290234 192402
rect 292110 192374 292138 192402
rect 292110 189854 292138 189882
rect 282646 149534 282674 149562
rect 288526 169694 288554 169722
rect 280966 72254 280994 72282
rect 297374 164206 297402 164234
rect 297374 163366 297402 163394
rect 297766 143262 297794 143290
rect 297766 113414 297794 113442
rect 290206 89894 290234 89922
rect 290206 81046 290234 81074
rect 297766 49966 297794 49994
rect 297878 29974 297906 30002
rect 297878 14798 297906 14826
rect 297766 14686 297794 14714
rect 288526 14070 288554 14098
rect 276766 9254 276794 9282
rect 257446 3374 257474 3402
<< metal3 >>
rect 15521 297878 15526 297906
rect 15554 297878 116662 297906
rect 116690 297878 116695 297906
rect 216561 297878 216566 297906
rect 216594 297878 255486 297906
rect 255514 297878 255519 297906
rect 32321 297822 32326 297850
rect 32354 297822 50134 297850
rect 50162 297822 50167 297850
rect 94593 297822 94598 297850
rect 94626 297822 221326 297850
rect 221354 297822 221359 297850
rect 275081 297822 275086 297850
rect 275114 297822 282982 297850
rect 283010 297822 283015 297850
rect 16361 297766 16366 297794
rect 16394 297766 294070 297794
rect 294098 297766 294103 297794
rect 299760 296548 300480 296660
rect 194385 295918 194390 295946
rect 194418 295918 196126 295946
rect 196154 295918 196159 295946
rect -480 295722 240 295820
rect -480 295708 2086 295722
rect 196 295694 2086 295708
rect 2114 295694 2119 295722
rect 183297 294406 183302 294434
rect 183330 294406 188566 294434
rect 188594 294406 188599 294434
rect 196121 291326 196126 291354
rect 196154 291326 199486 291354
rect 199514 291326 199519 291354
rect 299760 289898 300480 289996
rect 293986 289884 300480 289898
rect 293986 289870 299796 289884
rect 293986 289842 294014 289870
rect 10033 289814 10038 289842
rect 10066 289814 294014 289842
rect -480 288610 240 288708
rect -480 288596 5446 288610
rect 196 288582 5446 288596
rect 5474 288582 5479 288610
rect 80201 288526 80206 288554
rect 80234 288526 83174 288554
rect 83202 288526 83207 288554
rect 199481 287686 199486 287714
rect 199514 287686 201166 287714
rect 201194 287686 201199 287714
rect 188561 283878 188566 283906
rect 188594 283878 190246 283906
rect 190274 283878 190279 283906
rect 299760 283234 300480 283332
rect 293986 283220 300480 283234
rect 293986 283206 299796 283220
rect 293986 283122 294014 283206
rect 258281 283094 258286 283122
rect 258314 283094 294014 283122
rect 57129 281806 57134 281834
rect 57162 281806 80206 281834
rect 80234 281806 80239 281834
rect -480 281484 240 281596
rect 201161 280574 201166 280602
rect 201194 280574 204134 280602
rect 204162 280574 204167 280602
rect 52481 279286 52486 279314
rect 52514 279286 57134 279314
rect 57162 279286 57167 279314
rect 204129 278446 204134 278474
rect 204162 278446 206206 278474
rect 206234 278446 206239 278474
rect 299760 276556 300480 276668
rect 206201 275926 206206 275954
rect 206234 275926 219534 275954
rect 219562 275926 219567 275954
rect 23641 275086 23646 275114
rect 23674 275086 52486 275114
rect 52514 275086 52519 275114
rect -480 274386 240 274484
rect -480 274372 3766 274386
rect 196 274358 3766 274372
rect 3794 274358 3799 274386
rect 21009 272566 21014 272594
rect 21042 272566 23646 272594
rect 23674 272566 23679 272594
rect 219529 271726 219534 271754
rect 219562 271726 226366 271754
rect 226394 271726 226399 271754
rect 19721 271390 19726 271418
rect 19754 271390 21014 271418
rect 21042 271390 21047 271418
rect 299760 269906 300480 270004
rect 297761 269878 297766 269906
rect 297794 269892 300480 269906
rect 297794 269878 299796 269892
rect 190241 268366 190246 268394
rect 190274 268366 196966 268394
rect 196994 268366 196999 268394
rect 18489 267974 18494 268002
rect 18522 267974 19726 268002
rect 19754 267974 19759 268002
rect -480 267274 240 267372
rect -480 267260 5894 267274
rect 196 267246 5894 267260
rect 5866 267162 5894 267246
rect 5866 267134 7966 267162
rect 7994 267134 7999 267162
rect 17201 265846 17206 265874
rect 17234 265846 18438 265874
rect 18466 265846 18471 265874
rect 226361 265006 226366 265034
rect 226394 265006 233086 265034
rect 233114 265006 233119 265034
rect 299760 263242 300480 263340
rect 299726 263228 300480 263242
rect 299726 263214 299796 263228
rect 299726 263186 299754 263214
rect 299726 263158 299810 263186
rect 299782 262962 299810 263158
rect 282641 262934 282646 262962
rect 282674 262934 299810 262962
rect 233081 262486 233086 262514
rect 233114 262486 236614 262514
rect 236642 262486 236647 262514
rect 14625 261646 14630 261674
rect 14658 261646 17206 261674
rect 17234 261646 17239 261674
rect 236609 260358 236614 260386
rect 236642 260358 238966 260386
rect 238994 260358 238999 260386
rect -480 260148 240 260260
rect 10873 260022 10878 260050
rect 10906 260022 160454 260050
rect 160482 260022 160487 260050
rect 12553 259966 12558 259994
rect 12586 259966 260414 259994
rect 260442 259966 260447 259994
rect 16809 259182 16814 259210
rect 16842 259182 105854 259210
rect 105882 259182 105892 259210
rect 5441 259126 5446 259154
rect 5474 259126 180614 259154
rect 180642 259126 180647 259154
rect 196961 258454 196966 258482
rect 196994 258454 231798 258482
rect 231826 258454 231831 258482
rect 230393 258398 230398 258426
rect 230426 258398 282646 258426
rect 282674 258398 282679 258426
rect 14289 258342 14294 258370
rect 14322 258342 149534 258370
rect 149562 258342 149567 258370
rect 188729 258342 188734 258370
rect 188762 258342 258286 258370
rect 258314 258342 258319 258370
rect 13337 258286 13342 258314
rect 13370 258286 297766 258314
rect 297794 258286 297799 258314
rect 97673 257502 97678 257530
rect 97706 257502 226814 257530
rect 226842 257502 226847 257530
rect 231793 257502 231798 257530
rect 231826 257502 255150 257530
rect 255178 257502 255183 257530
rect 2081 257446 2086 257474
rect 2114 257446 257054 257474
rect 257082 257446 257087 257474
rect 221321 257110 221326 257138
rect 221354 257110 221774 257138
rect 221802 257110 221807 257138
rect 14681 257054 14686 257082
rect 14714 257054 255038 257082
rect 255066 257054 255071 257082
rect 31481 256718 31486 256746
rect 31514 256718 32326 256746
rect 32354 256718 32359 256746
rect 238961 256606 238966 256634
rect 238994 256606 254870 256634
rect 254898 256606 254903 256634
rect 23081 256550 23086 256578
rect 23114 256550 279286 256578
rect 279314 256550 279319 256578
rect 299760 256564 300480 256676
rect 155801 256494 155806 256522
rect 155834 256494 258286 256522
rect 258314 256494 258319 256522
rect 8913 256438 8918 256466
rect 8946 256438 163870 256466
rect 163898 256438 163903 256466
rect 197129 256438 197134 256466
rect 197162 256438 280126 256466
rect 280154 256438 280159 256466
rect 6281 256382 6286 256410
rect 6314 256382 213374 256410
rect 213402 256382 213407 256410
rect 39545 256326 39550 256354
rect 39578 256326 61670 256354
rect 61698 256326 61703 256354
rect 64409 256326 64414 256354
rect 64442 256326 282646 256354
rect 282674 256326 282679 256354
rect 7177 256270 7182 256298
rect 7210 256270 238070 256298
rect 238098 256270 238103 256298
rect 2193 255878 2198 255906
rect 2226 255878 130550 255906
rect 130578 255878 130583 255906
rect 249489 255878 249494 255906
rect 249522 255878 255374 255906
rect 255402 255878 255407 255906
rect 14457 255822 14462 255850
rect 14490 255822 27734 255850
rect 27762 255822 27767 255850
rect 127689 255822 127694 255850
rect 127722 255822 255430 255850
rect 255458 255822 255463 255850
rect 14345 255766 14350 255794
rect 14378 255766 60494 255794
rect 60522 255766 60527 255794
rect 61665 255766 61670 255794
rect 61698 255766 297766 255794
rect 297794 255766 297799 255794
rect 14177 255654 14182 255682
rect 14210 255654 16366 255682
rect 16394 255654 16399 255682
rect 172265 255542 172270 255570
rect 172298 255542 262486 255570
rect 262514 255542 262519 255570
rect 5441 255486 5446 255514
rect 5474 255486 122150 255514
rect 122178 255486 122183 255514
rect 147401 255486 147406 255514
rect 147434 255486 267526 255514
rect 267554 255486 267559 255514
rect 89273 255430 89278 255458
rect 89306 255430 266686 255458
rect 266714 255430 266719 255458
rect 15185 255374 15190 255402
rect 15218 255374 260862 255402
rect 260890 255374 260895 255402
rect 12497 255206 12502 255234
rect 12530 255206 17654 255234
rect 17626 255178 17654 255206
rect 13393 255150 13398 255178
rect 13426 255150 15526 255178
rect 15554 255150 15559 255178
rect 17626 255150 297822 255178
rect 297850 255150 297855 255178
rect 2137 255094 2142 255122
rect 2170 255094 257110 255122
rect 257138 255094 257143 255122
rect 14737 253638 14742 253666
rect 14770 253638 15190 253666
rect 15218 253638 15223 253666
rect -480 253050 240 253148
rect -480 253036 266 253050
rect 196 253022 266 253036
rect 238 252994 266 253022
rect 182 252966 266 252994
rect 182 252882 210 252966
rect 182 252854 7126 252882
rect 7154 252854 7159 252882
rect 14233 252014 14238 252042
rect 14266 252014 14686 252042
rect 14714 252014 14719 252042
rect 14121 251174 14126 251202
rect 14154 251174 14742 251202
rect 14770 251174 14775 251202
rect 299760 249914 300480 250012
rect 299726 249900 300480 249914
rect 299726 249886 299796 249900
rect 299726 249858 299754 249886
rect 299726 249830 299810 249858
rect 299782 249522 299810 249830
rect 260801 249494 260806 249522
rect 260834 249494 299810 249522
rect 260857 248206 260862 248234
rect 260890 248206 265846 248234
rect 265874 248206 265879 248234
rect 254884 246862 257446 246890
rect 257474 246862 257479 246890
rect 15134 246162 15162 246820
rect 8857 246134 8862 246162
rect 8890 246134 15162 246162
rect -480 245938 240 246036
rect -480 245924 266 245938
rect 196 245910 266 245924
rect 238 245882 266 245910
rect 182 245854 266 245882
rect 182 245322 210 245854
rect 2081 245686 2086 245714
rect 2114 245686 8918 245714
rect 8946 245686 8951 245714
rect 265841 245686 265846 245714
rect 265874 245686 270606 245714
rect 270634 245686 270639 245714
rect 182 245294 8806 245322
rect 8834 245294 8839 245322
rect 297817 243334 297822 243362
rect 297850 243348 299796 243362
rect 297850 243334 300480 243348
rect 299760 243236 300480 243334
rect 270601 243166 270606 243194
rect 270634 243166 279342 243194
rect 279370 243166 279375 243194
rect 279337 239806 279342 239834
rect 279370 239806 297822 239834
rect 297850 239806 297855 239834
rect -480 238812 240 238924
rect 254884 238462 257110 238490
rect 257138 238462 257143 238490
rect 15134 237762 15162 238420
rect 7121 237734 7126 237762
rect 7154 237734 15162 237762
rect 299760 236572 300480 236684
rect 196 231812 2198 231826
rect -480 231798 2198 231812
rect 2226 231798 2231 231826
rect -480 231700 240 231798
rect 14457 230398 14462 230426
rect 14490 230398 15148 230426
rect 254884 230398 258734 230426
rect 258706 230202 258734 230398
rect 258706 230174 259126 230202
rect 259154 230174 259159 230202
rect 297817 230006 297822 230034
rect 297850 230020 299796 230034
rect 297850 230006 300480 230020
rect 299760 229908 300480 230006
rect -480 224602 240 224700
rect -480 224588 2198 224602
rect 196 224574 2198 224588
rect 2226 224574 2231 224602
rect 255033 224238 255038 224266
rect 255066 224238 256606 224266
rect 256634 224238 256639 224266
rect 297761 223342 297766 223370
rect 297794 223356 299796 223370
rect 297794 223342 300480 223356
rect 299760 223244 300480 223342
rect 15134 221802 15162 221956
rect 5889 221774 5894 221802
rect 5922 221774 15162 221802
rect 256601 219646 256606 219674
rect 256634 219646 274246 219674
rect 274274 219646 274279 219674
rect -480 217476 240 217588
rect 299760 216580 300480 216692
rect 274241 212926 274246 212954
rect 274274 212926 280182 212954
rect 280210 212926 280215 212954
rect 196 210476 2142 210490
rect -480 210462 2142 210476
rect 2170 210462 2175 210490
rect -480 210364 240 210462
rect 299760 209930 300480 210028
rect 299726 209916 300480 209930
rect 299726 209902 299796 209916
rect 299726 209874 299754 209902
rect 299726 209846 299810 209874
rect 280177 209566 280182 209594
rect 280210 209566 284326 209594
rect 284354 209566 284359 209594
rect 299782 209202 299810 209846
rect 268361 209174 268366 209202
rect 268394 209174 299810 209202
rect 254884 205534 255486 205562
rect 255514 205534 255519 205562
rect -480 203322 240 203364
rect 299760 203322 300480 203364
rect -480 203294 6286 203322
rect 6314 203294 6319 203322
rect 280961 203294 280966 203322
rect 280994 203294 300480 203322
rect -480 203252 240 203294
rect 299760 203252 300480 203294
rect 284321 200718 284326 200746
rect 284354 200718 286846 200746
rect 286874 200718 286879 200746
rect 15134 196602 15162 197092
rect 7121 196574 7126 196602
rect 7154 196574 15162 196602
rect 299760 196588 300480 196700
rect -480 196140 240 196252
rect 286841 194446 286846 194474
rect 286874 194446 290206 194474
rect 290234 194446 290239 194474
rect 290201 192374 290206 192402
rect 290234 192374 292110 192402
rect 292138 192374 292143 192402
rect 299760 189938 300480 190036
rect 293986 189924 300480 189938
rect 293986 189910 299796 189924
rect 293986 189882 294014 189910
rect 292105 189854 292110 189882
rect 292138 189854 294014 189882
rect -480 189042 240 189140
rect -480 189028 3822 189042
rect 196 189014 3822 189028
rect 3850 189014 3855 189042
rect 14121 188734 14126 188762
rect 14154 188734 15148 188762
rect 254884 188734 258734 188762
rect 258706 188202 258734 188734
rect 258706 188174 275086 188202
rect 275114 188174 275119 188202
rect 299760 183274 300480 183372
rect 293986 183260 300480 183274
rect 293986 183246 299796 183260
rect 293986 183162 294014 183246
rect 262481 183134 262486 183162
rect 262514 183134 294014 183162
rect 196 182028 2086 182042
rect -480 182014 2086 182028
rect 2114 182014 2119 182042
rect -480 181916 240 182014
rect 14345 180670 14350 180698
rect 14378 180670 15148 180698
rect 299760 176596 300480 176708
rect -480 174804 240 174916
rect 299760 169946 300480 170044
rect 299726 169932 300480 169946
rect 299726 169918 299796 169932
rect 299726 169890 299754 169918
rect 299726 169862 299810 169890
rect 299782 169722 299810 169862
rect 288521 169694 288526 169722
rect 288554 169694 299810 169722
rect 196 167804 5446 167818
rect -480 167790 5446 167804
rect 5474 167790 5479 167818
rect -480 167692 240 167790
rect 258281 164206 258286 164234
rect 258314 164206 297374 164234
rect 297402 164206 297407 164234
rect 14177 163870 14182 163898
rect 14210 163870 15148 163898
rect 254884 163870 257894 163898
rect 257922 163870 257927 163898
rect 297369 163366 297374 163394
rect 297402 163380 299796 163394
rect 297402 163366 300480 163380
rect 299760 163268 300480 163366
rect -480 160594 240 160692
rect -480 160580 5894 160594
rect 196 160566 5894 160580
rect 5866 160482 5894 160566
rect 5866 160454 7182 160482
rect 7210 160454 7215 160482
rect 299760 156604 300480 156716
rect 15134 155442 15162 155764
rect 5497 155414 5502 155442
rect 5530 155414 15162 155442
rect -480 153468 240 153580
rect 299760 149954 300480 150052
rect 299726 149940 300480 149954
rect 299726 149926 299796 149940
rect 299726 149898 299754 149926
rect 299726 149870 299810 149898
rect 299782 149562 299810 149870
rect 282641 149534 282646 149562
rect 282674 149534 299810 149562
rect 12497 147406 12502 147434
rect 12530 147406 15148 147434
rect 254884 147406 258286 147434
rect 258314 147406 258319 147434
rect -480 146370 240 146468
rect -480 146356 5446 146370
rect 196 146342 5446 146356
rect 5474 146342 5479 146370
rect 299760 143290 300480 143388
rect 297761 143262 297766 143290
rect 297794 143276 300480 143290
rect 297794 143262 299796 143276
rect -480 139258 240 139356
rect -480 139244 2086 139258
rect 196 139230 2086 139244
rect 2114 139230 2119 139258
rect 2193 139006 2198 139034
rect 2226 139006 8022 139034
rect 8050 139006 8055 139034
rect 13337 139006 13342 139034
rect 13370 139006 15148 139034
rect 254884 139006 255766 139034
rect 255794 139006 255799 139034
rect 299760 136612 300480 136724
rect -480 132132 240 132244
rect 254884 130942 257110 130970
rect 257138 130942 257143 130970
rect 299760 129962 300480 130060
rect 299726 129948 300480 129962
rect 299726 129934 299796 129948
rect 299726 129906 299754 129934
rect 299726 129878 299810 129906
rect 299782 129402 299810 129878
rect 279281 129374 279286 129402
rect 279314 129374 299810 129402
rect -480 125034 240 125132
rect -480 125020 2142 125034
rect 196 125006 2142 125020
rect 2170 125006 2175 125034
rect 299760 123298 300480 123396
rect 299726 123284 300480 123298
rect 299726 123270 299796 123284
rect 299726 123242 299754 123270
rect 299726 123214 299810 123242
rect 299782 122682 299810 123214
rect 267521 122654 267526 122682
rect 267554 122654 299810 122682
rect 254884 122542 257054 122570
rect 257082 122542 257087 122570
rect -480 117922 240 118020
rect -480 117908 266 117922
rect 196 117894 266 117908
rect 238 117866 266 117894
rect 182 117838 266 117866
rect 182 117642 210 117838
rect 182 117614 8862 117642
rect 8890 117614 8895 117642
rect 299760 116620 300480 116732
rect 254884 114142 256662 114170
rect 256690 114142 256695 114170
rect 256657 113414 256662 113442
rect 256690 113414 297766 113442
rect 297794 113414 297799 113442
rect -480 110796 240 110908
rect 299760 109970 300480 110068
rect 299726 109956 300480 109970
rect 299726 109942 299796 109956
rect 299726 109914 299754 109942
rect 299726 109886 299810 109914
rect 299782 109242 299810 109886
rect 280121 109214 280126 109242
rect 280154 109214 299810 109242
rect 254884 106078 258734 106106
rect 14345 106022 14350 106050
rect 14378 106022 15148 106050
rect 258706 105882 258734 106078
rect 258706 105854 276766 105882
rect 276794 105854 276799 105882
rect 196 103796 5502 103810
rect -480 103782 5502 103796
rect 5530 103782 5535 103810
rect -480 103684 240 103782
rect 299760 103362 300480 103404
rect 258281 103334 258286 103362
rect 258314 103334 300480 103362
rect 299760 103292 300480 103334
rect 254884 97678 258734 97706
rect 13449 97622 13454 97650
rect 13482 97622 15148 97650
rect 258706 97482 258734 97678
rect 258706 97454 261646 97482
rect 261674 97454 261679 97482
rect -480 96642 240 96684
rect -480 96614 13454 96642
rect 13482 96614 13487 96642
rect 299760 96628 300480 96740
rect -480 96572 240 96614
rect 299760 89978 300480 90076
rect 293986 89964 300480 89978
rect 293986 89950 299796 89964
rect 293986 89922 294014 89950
rect 290201 89894 290206 89922
rect 290234 89894 294014 89922
rect -480 89460 240 89572
rect 254884 89278 258286 89306
rect 258314 89278 258319 89306
rect 12161 89222 12166 89250
rect 12194 89222 15148 89250
rect 299760 83314 300480 83412
rect 293986 83300 300480 83314
rect 293986 83286 299796 83300
rect 293986 83202 294014 83286
rect 261641 83174 261646 83202
rect 261674 83174 294014 83202
rect -480 82362 240 82460
rect -480 82348 14686 82362
rect 196 82334 14686 82348
rect 14714 82334 14719 82362
rect 14233 81214 14238 81242
rect 14266 81214 15148 81242
rect 280569 81046 280574 81074
rect 280602 81046 290206 81074
rect 290234 81046 290239 81074
rect 275921 77686 275926 77714
rect 275954 77686 280574 77714
rect 280602 77686 280607 77714
rect 299760 76636 300480 76748
rect -480 75250 240 75348
rect -480 75236 266 75250
rect 196 75222 266 75236
rect 238 75194 266 75222
rect 182 75166 266 75194
rect 182 74802 210 75166
rect 182 74774 10486 74802
rect 10514 74774 10519 74802
rect 254884 72814 258734 72842
rect 14233 72758 14238 72786
rect 14266 72758 15148 72786
rect 258706 72282 258734 72814
rect 258706 72254 280966 72282
rect 280994 72254 280999 72282
rect 299760 69986 300480 70084
rect 299726 69972 300480 69986
rect 299726 69958 299796 69972
rect 299726 69930 299754 69958
rect 299726 69902 299810 69930
rect 299782 69762 299810 69902
rect 261641 69734 261646 69762
rect 261674 69734 299810 69762
rect -480 68124 240 68236
rect 14289 64414 14294 64442
rect 14322 64414 15148 64442
rect 299760 63322 300480 63420
rect 299726 63308 300480 63322
rect 299726 63294 299796 63308
rect 299726 63266 299754 63294
rect 299726 63238 299810 63266
rect 299782 63042 299810 63238
rect 266681 63014 266686 63042
rect 266714 63014 299810 63042
rect -480 61026 240 61124
rect -480 61012 2310 61026
rect 196 60998 2310 61012
rect 2338 60998 2343 61026
rect 299760 56644 300480 56756
rect 12553 56350 12558 56378
rect 12586 56350 15148 56378
rect 254884 56350 258734 56378
rect 258706 56322 258734 56350
rect 258706 56294 260806 56322
rect 260834 56294 260839 56322
rect 2305 54166 2310 54194
rect 2338 54166 12222 54194
rect 12250 54166 12255 54194
rect -480 53914 240 54012
rect -480 53900 2198 53914
rect 196 53886 2198 53900
rect 2226 53886 2231 53914
rect 273737 51254 273742 51282
rect 273770 51254 275926 51282
rect 275954 51254 275959 51282
rect 299760 49994 300480 50092
rect 297761 49966 297766 49994
rect 297794 49980 300480 49994
rect 297794 49966 299796 49980
rect 271721 48678 271726 48706
rect 271754 48678 273742 48706
rect 273770 48678 273775 48706
rect 254884 47950 256214 47978
rect 256242 47950 256247 47978
rect 10873 47894 10878 47922
rect 10906 47894 15148 47922
rect -480 46788 240 46900
rect 299760 43330 300480 43428
rect 299726 43316 300480 43330
rect 299726 43302 299796 43316
rect 299726 43274 299754 43302
rect 299726 43246 299810 43274
rect 299782 42882 299810 43246
rect 258281 42854 258286 42882
rect 258314 42854 299810 42882
rect 255089 42742 255094 42770
rect 255122 42742 256214 42770
rect 256242 42742 256247 42770
rect 270041 42406 270046 42434
rect 270074 42406 271726 42434
rect 271754 42406 271759 42434
rect -480 39690 240 39788
rect -480 39676 2310 39690
rect 196 39662 2310 39676
rect 2338 39662 2343 39690
rect 254884 39550 254982 39578
rect 255010 39550 255015 39578
rect 3761 39494 3766 39522
rect 3794 39494 15148 39522
rect 265841 39494 265846 39522
rect 265874 39494 270046 39522
rect 270074 39494 270079 39522
rect 299760 36652 300480 36764
rect 2305 36078 2310 36106
rect 2338 36078 4606 36106
rect 4634 36078 4639 36106
rect 260801 34846 260806 34874
rect 260834 34846 265846 34874
rect 265874 34846 265879 34874
rect 4601 33110 4606 33138
rect 4634 33110 5054 33138
rect 5082 33110 5087 33138
rect -480 32578 240 32676
rect -480 32564 266 32578
rect 196 32550 266 32564
rect 238 32522 266 32550
rect 182 32494 266 32522
rect 182 31962 210 32494
rect 2081 32326 2086 32354
rect 2114 32326 2926 32354
rect 2954 32326 2959 32354
rect 182 31934 12166 31962
rect 12194 31934 12199 31962
rect 2137 31878 2142 31906
rect 2170 31878 3262 31906
rect 3290 31878 3295 31906
rect 15134 31122 15162 31444
rect 7961 31094 7966 31122
rect 7994 31094 15162 31122
rect 5049 30646 5054 30674
rect 5082 30646 6846 30674
rect 6874 30646 6879 30674
rect 6841 30030 6846 30058
rect 6874 30030 7966 30058
rect 7994 30030 7999 30058
rect 299760 30002 300480 30100
rect 297873 29974 297878 30002
rect 297906 29988 300480 30002
rect 297906 29974 299796 29988
rect 3257 29806 3262 29834
rect 3290 29806 6286 29834
rect 6314 29806 6319 29834
rect 256601 29806 256606 29834
rect 256634 29806 260806 29834
rect 260834 29806 260839 29834
rect 7961 27734 7966 27762
rect 7994 27734 8862 27762
rect 8890 27734 8895 27762
rect 6281 26894 6286 26922
rect 6314 26894 6762 26922
rect 6734 26866 6762 26894
rect 6734 26838 9254 26866
rect 9282 26838 9287 26866
rect 255033 25886 255038 25914
rect 255066 25886 256606 25914
rect 256634 25886 256639 25914
rect -480 25452 240 25564
rect 9249 25158 9254 25186
rect 9282 25158 10934 25186
rect 10962 25158 10967 25186
rect 2921 24318 2926 24346
rect 2954 24318 3766 24346
rect 3794 24318 3799 24346
rect 10929 23926 10934 23954
rect 10962 23926 13006 23954
rect 13034 23926 13039 23954
rect 299760 23338 300480 23436
rect 299726 23324 300480 23338
rect 299726 23310 299796 23324
rect 299726 23282 299754 23310
rect 299726 23254 299810 23282
rect 254884 23086 255430 23114
rect 255458 23086 255463 23114
rect 15134 22722 15162 23044
rect 299782 22722 299810 23254
rect 10033 22694 10038 22722
rect 10066 22694 15162 22722
rect 259121 22694 259126 22722
rect 259154 22694 299810 22722
rect 3761 21406 3766 21434
rect 3794 21406 6958 21434
rect 6986 21406 6991 21434
rect 13001 21014 13006 21042
rect 13034 21014 13902 21042
rect 13930 21014 13935 21042
rect 8857 20958 8862 20986
rect 8890 20958 10934 20986
rect 10962 20958 10967 20986
rect 10929 19726 10934 19754
rect 10962 19726 12166 19754
rect 12194 19726 12199 19754
rect 13897 19278 13902 19306
rect 13930 19278 14742 19306
rect 14770 19278 14775 19306
rect 12161 18494 12166 18522
rect 12194 18494 13482 18522
rect 13454 18466 13482 18494
rect -480 18354 240 18452
rect 13454 18438 14910 18466
rect 14938 18438 14943 18466
rect -480 18340 266 18354
rect 196 18326 266 18340
rect 238 18298 266 18326
rect 182 18270 266 18298
rect 182 17682 210 18270
rect 6953 18046 6958 18074
rect 6986 18046 14798 18074
rect 14826 18046 14831 18074
rect 182 17654 7126 17682
rect 7154 17654 7159 17682
rect 299760 16660 300480 16772
rect 13393 15918 13398 15946
rect 13426 15918 14966 15946
rect 14994 15918 14999 15946
rect 2193 15526 2198 15554
rect 2226 15526 15274 15554
rect 15246 15106 15274 15526
rect 15241 15078 15246 15106
rect 15274 15078 15279 15106
rect 14793 14910 14798 14938
rect 14826 14910 255094 14938
rect 255122 14910 255127 14938
rect 14905 14854 14910 14882
rect 14938 14854 254982 14882
rect 255010 14854 255015 14882
rect 14345 14798 14350 14826
rect 14378 14798 297878 14826
rect 297906 14798 297911 14826
rect 166105 14686 166110 14714
rect 166138 14686 297766 14714
rect 297794 14686 297799 14714
rect 10481 14462 10486 14490
rect 10514 14462 64358 14490
rect 64386 14462 64391 14490
rect 14681 14406 14686 14434
rect 14714 14406 72758 14434
rect 72786 14406 72791 14434
rect 5441 14350 5446 14378
rect 5474 14350 163814 14378
rect 163842 14350 163847 14378
rect 197129 14350 197134 14378
rect 197162 14350 268366 14378
rect 268394 14350 268399 14378
rect 3817 14294 3822 14322
rect 3850 14294 246806 14322
rect 246834 14294 246839 14322
rect 8017 14238 8022 14266
rect 8050 14238 23030 14266
rect 23058 14238 23063 14266
rect 8801 14182 8806 14210
rect 8834 14182 56294 14210
rect 56322 14182 56327 14210
rect 81209 14182 81214 14210
rect 81242 14182 254870 14210
rect 254898 14182 254903 14210
rect 12217 14126 12222 14154
rect 12250 14126 106022 14154
rect 106050 14126 106055 14154
rect 147401 14126 147406 14154
rect 147434 14126 261646 14154
rect 261674 14126 261679 14154
rect 15241 14070 15246 14098
rect 15274 14070 97622 14098
rect 97650 14070 97655 14098
rect 130937 14070 130942 14098
rect 130970 14070 166110 14098
rect 166138 14070 166143 14098
rect 180665 14070 180670 14098
rect 180698 14070 288526 14098
rect 288554 14070 288559 14098
rect 221993 14014 221998 14042
rect 222026 14014 255374 14042
rect 255402 14014 255407 14042
rect 14289 13958 14294 13986
rect 14322 13958 255038 13986
rect 255066 13958 255071 13986
rect 7569 13846 7574 13874
rect 7602 13846 257110 13874
rect 257138 13846 257143 13874
rect 14737 13398 14742 13426
rect 14770 13398 255766 13426
rect 255794 13398 255799 13426
rect 14625 13342 14630 13370
rect 14658 13342 172214 13370
rect 172242 13342 172247 13370
rect 139001 13286 139006 13314
rect 139034 13286 255150 13314
rect 255178 13286 255183 13314
rect -480 11242 240 11340
rect -480 11228 266 11242
rect 196 11214 266 11228
rect 238 11186 266 11214
rect 182 11158 266 11186
rect 182 10962 210 11158
rect 182 10934 257894 10962
rect 257922 10934 257927 10962
rect 299760 10010 300480 10108
rect 299726 9996 300480 10010
rect 299726 9982 299796 9996
rect 299726 9954 299754 9982
rect 299726 9926 299810 9954
rect 299782 9282 299810 9926
rect 276761 9254 276766 9282
rect 276794 9254 299810 9282
rect -480 4116 240 4228
rect 299760 3402 300480 3444
rect 257441 3374 257446 3402
rect 257474 3374 300480 3402
rect 299760 3332 300480 3374
<< via3 >>
rect 254870 256606 254898 256634
rect 15190 255374 15218 255402
rect 15190 253638 15218 253666
rect 254870 14182 254898 14210
<< metal4 >>
rect -6 299670 304 299718
rect -6 299642 42 299670
rect 70 299642 104 299670
rect 132 299642 166 299670
rect 194 299642 228 299670
rect 256 299642 304 299670
rect -6 299608 304 299642
rect -6 299580 42 299608
rect 70 299580 104 299608
rect 132 299580 166 299608
rect 194 299580 228 299608
rect 256 299580 304 299608
rect -6 299546 304 299580
rect -6 299518 42 299546
rect 70 299518 104 299546
rect 132 299518 166 299546
rect 194 299518 228 299546
rect 256 299518 304 299546
rect -6 299484 304 299518
rect -6 299456 42 299484
rect 70 299456 104 299484
rect 132 299456 166 299484
rect 194 299456 228 299484
rect 256 299456 304 299484
rect -6 293959 304 299456
rect -6 293931 42 293959
rect 70 293931 104 293959
rect 132 293931 166 293959
rect 194 293931 228 293959
rect 256 293931 304 293959
rect -6 293897 304 293931
rect -6 293869 42 293897
rect 70 293869 104 293897
rect 132 293869 166 293897
rect 194 293869 228 293897
rect 256 293869 304 293897
rect -6 293835 304 293869
rect -6 293807 42 293835
rect 70 293807 104 293835
rect 132 293807 166 293835
rect 194 293807 228 293835
rect 256 293807 304 293835
rect -6 293773 304 293807
rect -6 293745 42 293773
rect 70 293745 104 293773
rect 132 293745 166 293773
rect 194 293745 228 293773
rect 256 293745 304 293773
rect -6 284959 304 293745
rect -6 284931 42 284959
rect 70 284931 104 284959
rect 132 284931 166 284959
rect 194 284931 228 284959
rect 256 284931 304 284959
rect -6 284897 304 284931
rect -6 284869 42 284897
rect 70 284869 104 284897
rect 132 284869 166 284897
rect 194 284869 228 284897
rect 256 284869 304 284897
rect -6 284835 304 284869
rect -6 284807 42 284835
rect 70 284807 104 284835
rect 132 284807 166 284835
rect 194 284807 228 284835
rect 256 284807 304 284835
rect -6 284773 304 284807
rect -6 284745 42 284773
rect 70 284745 104 284773
rect 132 284745 166 284773
rect 194 284745 228 284773
rect 256 284745 304 284773
rect -6 275959 304 284745
rect -6 275931 42 275959
rect 70 275931 104 275959
rect 132 275931 166 275959
rect 194 275931 228 275959
rect 256 275931 304 275959
rect -6 275897 304 275931
rect -6 275869 42 275897
rect 70 275869 104 275897
rect 132 275869 166 275897
rect 194 275869 228 275897
rect 256 275869 304 275897
rect -6 275835 304 275869
rect -6 275807 42 275835
rect 70 275807 104 275835
rect 132 275807 166 275835
rect 194 275807 228 275835
rect 256 275807 304 275835
rect -6 275773 304 275807
rect -6 275745 42 275773
rect 70 275745 104 275773
rect 132 275745 166 275773
rect 194 275745 228 275773
rect 256 275745 304 275773
rect -6 266959 304 275745
rect -6 266931 42 266959
rect 70 266931 104 266959
rect 132 266931 166 266959
rect 194 266931 228 266959
rect 256 266931 304 266959
rect -6 266897 304 266931
rect -6 266869 42 266897
rect 70 266869 104 266897
rect 132 266869 166 266897
rect 194 266869 228 266897
rect 256 266869 304 266897
rect -6 266835 304 266869
rect -6 266807 42 266835
rect 70 266807 104 266835
rect 132 266807 166 266835
rect 194 266807 228 266835
rect 256 266807 304 266835
rect -6 266773 304 266807
rect -6 266745 42 266773
rect 70 266745 104 266773
rect 132 266745 166 266773
rect 194 266745 228 266773
rect 256 266745 304 266773
rect -6 257959 304 266745
rect -6 257931 42 257959
rect 70 257931 104 257959
rect 132 257931 166 257959
rect 194 257931 228 257959
rect 256 257931 304 257959
rect -6 257897 304 257931
rect -6 257869 42 257897
rect 70 257869 104 257897
rect 132 257869 166 257897
rect 194 257869 228 257897
rect 256 257869 304 257897
rect -6 257835 304 257869
rect -6 257807 42 257835
rect 70 257807 104 257835
rect 132 257807 166 257835
rect 194 257807 228 257835
rect 256 257807 304 257835
rect -6 257773 304 257807
rect -6 257745 42 257773
rect 70 257745 104 257773
rect 132 257745 166 257773
rect 194 257745 228 257773
rect 256 257745 304 257773
rect -6 248959 304 257745
rect -6 248931 42 248959
rect 70 248931 104 248959
rect 132 248931 166 248959
rect 194 248931 228 248959
rect 256 248931 304 248959
rect -6 248897 304 248931
rect -6 248869 42 248897
rect 70 248869 104 248897
rect 132 248869 166 248897
rect 194 248869 228 248897
rect 256 248869 304 248897
rect -6 248835 304 248869
rect -6 248807 42 248835
rect 70 248807 104 248835
rect 132 248807 166 248835
rect 194 248807 228 248835
rect 256 248807 304 248835
rect -6 248773 304 248807
rect -6 248745 42 248773
rect 70 248745 104 248773
rect 132 248745 166 248773
rect 194 248745 228 248773
rect 256 248745 304 248773
rect -6 239959 304 248745
rect -6 239931 42 239959
rect 70 239931 104 239959
rect 132 239931 166 239959
rect 194 239931 228 239959
rect 256 239931 304 239959
rect -6 239897 304 239931
rect -6 239869 42 239897
rect 70 239869 104 239897
rect 132 239869 166 239897
rect 194 239869 228 239897
rect 256 239869 304 239897
rect -6 239835 304 239869
rect -6 239807 42 239835
rect 70 239807 104 239835
rect 132 239807 166 239835
rect 194 239807 228 239835
rect 256 239807 304 239835
rect -6 239773 304 239807
rect -6 239745 42 239773
rect 70 239745 104 239773
rect 132 239745 166 239773
rect 194 239745 228 239773
rect 256 239745 304 239773
rect -6 230959 304 239745
rect -6 230931 42 230959
rect 70 230931 104 230959
rect 132 230931 166 230959
rect 194 230931 228 230959
rect 256 230931 304 230959
rect -6 230897 304 230931
rect -6 230869 42 230897
rect 70 230869 104 230897
rect 132 230869 166 230897
rect 194 230869 228 230897
rect 256 230869 304 230897
rect -6 230835 304 230869
rect -6 230807 42 230835
rect 70 230807 104 230835
rect 132 230807 166 230835
rect 194 230807 228 230835
rect 256 230807 304 230835
rect -6 230773 304 230807
rect -6 230745 42 230773
rect 70 230745 104 230773
rect 132 230745 166 230773
rect 194 230745 228 230773
rect 256 230745 304 230773
rect -6 221959 304 230745
rect -6 221931 42 221959
rect 70 221931 104 221959
rect 132 221931 166 221959
rect 194 221931 228 221959
rect 256 221931 304 221959
rect -6 221897 304 221931
rect -6 221869 42 221897
rect 70 221869 104 221897
rect 132 221869 166 221897
rect 194 221869 228 221897
rect 256 221869 304 221897
rect -6 221835 304 221869
rect -6 221807 42 221835
rect 70 221807 104 221835
rect 132 221807 166 221835
rect 194 221807 228 221835
rect 256 221807 304 221835
rect -6 221773 304 221807
rect -6 221745 42 221773
rect 70 221745 104 221773
rect 132 221745 166 221773
rect 194 221745 228 221773
rect 256 221745 304 221773
rect -6 212959 304 221745
rect -6 212931 42 212959
rect 70 212931 104 212959
rect 132 212931 166 212959
rect 194 212931 228 212959
rect 256 212931 304 212959
rect -6 212897 304 212931
rect -6 212869 42 212897
rect 70 212869 104 212897
rect 132 212869 166 212897
rect 194 212869 228 212897
rect 256 212869 304 212897
rect -6 212835 304 212869
rect -6 212807 42 212835
rect 70 212807 104 212835
rect 132 212807 166 212835
rect 194 212807 228 212835
rect 256 212807 304 212835
rect -6 212773 304 212807
rect -6 212745 42 212773
rect 70 212745 104 212773
rect 132 212745 166 212773
rect 194 212745 228 212773
rect 256 212745 304 212773
rect -6 203959 304 212745
rect -6 203931 42 203959
rect 70 203931 104 203959
rect 132 203931 166 203959
rect 194 203931 228 203959
rect 256 203931 304 203959
rect -6 203897 304 203931
rect -6 203869 42 203897
rect 70 203869 104 203897
rect 132 203869 166 203897
rect 194 203869 228 203897
rect 256 203869 304 203897
rect -6 203835 304 203869
rect -6 203807 42 203835
rect 70 203807 104 203835
rect 132 203807 166 203835
rect 194 203807 228 203835
rect 256 203807 304 203835
rect -6 203773 304 203807
rect -6 203745 42 203773
rect 70 203745 104 203773
rect 132 203745 166 203773
rect 194 203745 228 203773
rect 256 203745 304 203773
rect -6 194959 304 203745
rect -6 194931 42 194959
rect 70 194931 104 194959
rect 132 194931 166 194959
rect 194 194931 228 194959
rect 256 194931 304 194959
rect -6 194897 304 194931
rect -6 194869 42 194897
rect 70 194869 104 194897
rect 132 194869 166 194897
rect 194 194869 228 194897
rect 256 194869 304 194897
rect -6 194835 304 194869
rect -6 194807 42 194835
rect 70 194807 104 194835
rect 132 194807 166 194835
rect 194 194807 228 194835
rect 256 194807 304 194835
rect -6 194773 304 194807
rect -6 194745 42 194773
rect 70 194745 104 194773
rect 132 194745 166 194773
rect 194 194745 228 194773
rect 256 194745 304 194773
rect -6 185959 304 194745
rect -6 185931 42 185959
rect 70 185931 104 185959
rect 132 185931 166 185959
rect 194 185931 228 185959
rect 256 185931 304 185959
rect -6 185897 304 185931
rect -6 185869 42 185897
rect 70 185869 104 185897
rect 132 185869 166 185897
rect 194 185869 228 185897
rect 256 185869 304 185897
rect -6 185835 304 185869
rect -6 185807 42 185835
rect 70 185807 104 185835
rect 132 185807 166 185835
rect 194 185807 228 185835
rect 256 185807 304 185835
rect -6 185773 304 185807
rect -6 185745 42 185773
rect 70 185745 104 185773
rect 132 185745 166 185773
rect 194 185745 228 185773
rect 256 185745 304 185773
rect -6 176959 304 185745
rect -6 176931 42 176959
rect 70 176931 104 176959
rect 132 176931 166 176959
rect 194 176931 228 176959
rect 256 176931 304 176959
rect -6 176897 304 176931
rect -6 176869 42 176897
rect 70 176869 104 176897
rect 132 176869 166 176897
rect 194 176869 228 176897
rect 256 176869 304 176897
rect -6 176835 304 176869
rect -6 176807 42 176835
rect 70 176807 104 176835
rect 132 176807 166 176835
rect 194 176807 228 176835
rect 256 176807 304 176835
rect -6 176773 304 176807
rect -6 176745 42 176773
rect 70 176745 104 176773
rect 132 176745 166 176773
rect 194 176745 228 176773
rect 256 176745 304 176773
rect -6 167959 304 176745
rect -6 167931 42 167959
rect 70 167931 104 167959
rect 132 167931 166 167959
rect 194 167931 228 167959
rect 256 167931 304 167959
rect -6 167897 304 167931
rect -6 167869 42 167897
rect 70 167869 104 167897
rect 132 167869 166 167897
rect 194 167869 228 167897
rect 256 167869 304 167897
rect -6 167835 304 167869
rect -6 167807 42 167835
rect 70 167807 104 167835
rect 132 167807 166 167835
rect 194 167807 228 167835
rect 256 167807 304 167835
rect -6 167773 304 167807
rect -6 167745 42 167773
rect 70 167745 104 167773
rect 132 167745 166 167773
rect 194 167745 228 167773
rect 256 167745 304 167773
rect -6 158959 304 167745
rect -6 158931 42 158959
rect 70 158931 104 158959
rect 132 158931 166 158959
rect 194 158931 228 158959
rect 256 158931 304 158959
rect -6 158897 304 158931
rect -6 158869 42 158897
rect 70 158869 104 158897
rect 132 158869 166 158897
rect 194 158869 228 158897
rect 256 158869 304 158897
rect -6 158835 304 158869
rect -6 158807 42 158835
rect 70 158807 104 158835
rect 132 158807 166 158835
rect 194 158807 228 158835
rect 256 158807 304 158835
rect -6 158773 304 158807
rect -6 158745 42 158773
rect 70 158745 104 158773
rect 132 158745 166 158773
rect 194 158745 228 158773
rect 256 158745 304 158773
rect -6 149959 304 158745
rect -6 149931 42 149959
rect 70 149931 104 149959
rect 132 149931 166 149959
rect 194 149931 228 149959
rect 256 149931 304 149959
rect -6 149897 304 149931
rect -6 149869 42 149897
rect 70 149869 104 149897
rect 132 149869 166 149897
rect 194 149869 228 149897
rect 256 149869 304 149897
rect -6 149835 304 149869
rect -6 149807 42 149835
rect 70 149807 104 149835
rect 132 149807 166 149835
rect 194 149807 228 149835
rect 256 149807 304 149835
rect -6 149773 304 149807
rect -6 149745 42 149773
rect 70 149745 104 149773
rect 132 149745 166 149773
rect 194 149745 228 149773
rect 256 149745 304 149773
rect -6 140959 304 149745
rect -6 140931 42 140959
rect 70 140931 104 140959
rect 132 140931 166 140959
rect 194 140931 228 140959
rect 256 140931 304 140959
rect -6 140897 304 140931
rect -6 140869 42 140897
rect 70 140869 104 140897
rect 132 140869 166 140897
rect 194 140869 228 140897
rect 256 140869 304 140897
rect -6 140835 304 140869
rect -6 140807 42 140835
rect 70 140807 104 140835
rect 132 140807 166 140835
rect 194 140807 228 140835
rect 256 140807 304 140835
rect -6 140773 304 140807
rect -6 140745 42 140773
rect 70 140745 104 140773
rect 132 140745 166 140773
rect 194 140745 228 140773
rect 256 140745 304 140773
rect -6 131959 304 140745
rect -6 131931 42 131959
rect 70 131931 104 131959
rect 132 131931 166 131959
rect 194 131931 228 131959
rect 256 131931 304 131959
rect -6 131897 304 131931
rect -6 131869 42 131897
rect 70 131869 104 131897
rect 132 131869 166 131897
rect 194 131869 228 131897
rect 256 131869 304 131897
rect -6 131835 304 131869
rect -6 131807 42 131835
rect 70 131807 104 131835
rect 132 131807 166 131835
rect 194 131807 228 131835
rect 256 131807 304 131835
rect -6 131773 304 131807
rect -6 131745 42 131773
rect 70 131745 104 131773
rect 132 131745 166 131773
rect 194 131745 228 131773
rect 256 131745 304 131773
rect -6 122959 304 131745
rect -6 122931 42 122959
rect 70 122931 104 122959
rect 132 122931 166 122959
rect 194 122931 228 122959
rect 256 122931 304 122959
rect -6 122897 304 122931
rect -6 122869 42 122897
rect 70 122869 104 122897
rect 132 122869 166 122897
rect 194 122869 228 122897
rect 256 122869 304 122897
rect -6 122835 304 122869
rect -6 122807 42 122835
rect 70 122807 104 122835
rect 132 122807 166 122835
rect 194 122807 228 122835
rect 256 122807 304 122835
rect -6 122773 304 122807
rect -6 122745 42 122773
rect 70 122745 104 122773
rect 132 122745 166 122773
rect 194 122745 228 122773
rect 256 122745 304 122773
rect -6 113959 304 122745
rect -6 113931 42 113959
rect 70 113931 104 113959
rect 132 113931 166 113959
rect 194 113931 228 113959
rect 256 113931 304 113959
rect -6 113897 304 113931
rect -6 113869 42 113897
rect 70 113869 104 113897
rect 132 113869 166 113897
rect 194 113869 228 113897
rect 256 113869 304 113897
rect -6 113835 304 113869
rect -6 113807 42 113835
rect 70 113807 104 113835
rect 132 113807 166 113835
rect 194 113807 228 113835
rect 256 113807 304 113835
rect -6 113773 304 113807
rect -6 113745 42 113773
rect 70 113745 104 113773
rect 132 113745 166 113773
rect 194 113745 228 113773
rect 256 113745 304 113773
rect -6 104959 304 113745
rect -6 104931 42 104959
rect 70 104931 104 104959
rect 132 104931 166 104959
rect 194 104931 228 104959
rect 256 104931 304 104959
rect -6 104897 304 104931
rect -6 104869 42 104897
rect 70 104869 104 104897
rect 132 104869 166 104897
rect 194 104869 228 104897
rect 256 104869 304 104897
rect -6 104835 304 104869
rect -6 104807 42 104835
rect 70 104807 104 104835
rect 132 104807 166 104835
rect 194 104807 228 104835
rect 256 104807 304 104835
rect -6 104773 304 104807
rect -6 104745 42 104773
rect 70 104745 104 104773
rect 132 104745 166 104773
rect 194 104745 228 104773
rect 256 104745 304 104773
rect -6 95959 304 104745
rect -6 95931 42 95959
rect 70 95931 104 95959
rect 132 95931 166 95959
rect 194 95931 228 95959
rect 256 95931 304 95959
rect -6 95897 304 95931
rect -6 95869 42 95897
rect 70 95869 104 95897
rect 132 95869 166 95897
rect 194 95869 228 95897
rect 256 95869 304 95897
rect -6 95835 304 95869
rect -6 95807 42 95835
rect 70 95807 104 95835
rect 132 95807 166 95835
rect 194 95807 228 95835
rect 256 95807 304 95835
rect -6 95773 304 95807
rect -6 95745 42 95773
rect 70 95745 104 95773
rect 132 95745 166 95773
rect 194 95745 228 95773
rect 256 95745 304 95773
rect -6 86959 304 95745
rect -6 86931 42 86959
rect 70 86931 104 86959
rect 132 86931 166 86959
rect 194 86931 228 86959
rect 256 86931 304 86959
rect -6 86897 304 86931
rect -6 86869 42 86897
rect 70 86869 104 86897
rect 132 86869 166 86897
rect 194 86869 228 86897
rect 256 86869 304 86897
rect -6 86835 304 86869
rect -6 86807 42 86835
rect 70 86807 104 86835
rect 132 86807 166 86835
rect 194 86807 228 86835
rect 256 86807 304 86835
rect -6 86773 304 86807
rect -6 86745 42 86773
rect 70 86745 104 86773
rect 132 86745 166 86773
rect 194 86745 228 86773
rect 256 86745 304 86773
rect -6 77959 304 86745
rect -6 77931 42 77959
rect 70 77931 104 77959
rect 132 77931 166 77959
rect 194 77931 228 77959
rect 256 77931 304 77959
rect -6 77897 304 77931
rect -6 77869 42 77897
rect 70 77869 104 77897
rect 132 77869 166 77897
rect 194 77869 228 77897
rect 256 77869 304 77897
rect -6 77835 304 77869
rect -6 77807 42 77835
rect 70 77807 104 77835
rect 132 77807 166 77835
rect 194 77807 228 77835
rect 256 77807 304 77835
rect -6 77773 304 77807
rect -6 77745 42 77773
rect 70 77745 104 77773
rect 132 77745 166 77773
rect 194 77745 228 77773
rect 256 77745 304 77773
rect -6 68959 304 77745
rect -6 68931 42 68959
rect 70 68931 104 68959
rect 132 68931 166 68959
rect 194 68931 228 68959
rect 256 68931 304 68959
rect -6 68897 304 68931
rect -6 68869 42 68897
rect 70 68869 104 68897
rect 132 68869 166 68897
rect 194 68869 228 68897
rect 256 68869 304 68897
rect -6 68835 304 68869
rect -6 68807 42 68835
rect 70 68807 104 68835
rect 132 68807 166 68835
rect 194 68807 228 68835
rect 256 68807 304 68835
rect -6 68773 304 68807
rect -6 68745 42 68773
rect 70 68745 104 68773
rect 132 68745 166 68773
rect 194 68745 228 68773
rect 256 68745 304 68773
rect -6 59959 304 68745
rect -6 59931 42 59959
rect 70 59931 104 59959
rect 132 59931 166 59959
rect 194 59931 228 59959
rect 256 59931 304 59959
rect -6 59897 304 59931
rect -6 59869 42 59897
rect 70 59869 104 59897
rect 132 59869 166 59897
rect 194 59869 228 59897
rect 256 59869 304 59897
rect -6 59835 304 59869
rect -6 59807 42 59835
rect 70 59807 104 59835
rect 132 59807 166 59835
rect 194 59807 228 59835
rect 256 59807 304 59835
rect -6 59773 304 59807
rect -6 59745 42 59773
rect 70 59745 104 59773
rect 132 59745 166 59773
rect 194 59745 228 59773
rect 256 59745 304 59773
rect -6 50959 304 59745
rect -6 50931 42 50959
rect 70 50931 104 50959
rect 132 50931 166 50959
rect 194 50931 228 50959
rect 256 50931 304 50959
rect -6 50897 304 50931
rect -6 50869 42 50897
rect 70 50869 104 50897
rect 132 50869 166 50897
rect 194 50869 228 50897
rect 256 50869 304 50897
rect -6 50835 304 50869
rect -6 50807 42 50835
rect 70 50807 104 50835
rect 132 50807 166 50835
rect 194 50807 228 50835
rect 256 50807 304 50835
rect -6 50773 304 50807
rect -6 50745 42 50773
rect 70 50745 104 50773
rect 132 50745 166 50773
rect 194 50745 228 50773
rect 256 50745 304 50773
rect -6 41959 304 50745
rect -6 41931 42 41959
rect 70 41931 104 41959
rect 132 41931 166 41959
rect 194 41931 228 41959
rect 256 41931 304 41959
rect -6 41897 304 41931
rect -6 41869 42 41897
rect 70 41869 104 41897
rect 132 41869 166 41897
rect 194 41869 228 41897
rect 256 41869 304 41897
rect -6 41835 304 41869
rect -6 41807 42 41835
rect 70 41807 104 41835
rect 132 41807 166 41835
rect 194 41807 228 41835
rect 256 41807 304 41835
rect -6 41773 304 41807
rect -6 41745 42 41773
rect 70 41745 104 41773
rect 132 41745 166 41773
rect 194 41745 228 41773
rect 256 41745 304 41773
rect -6 32959 304 41745
rect -6 32931 42 32959
rect 70 32931 104 32959
rect 132 32931 166 32959
rect 194 32931 228 32959
rect 256 32931 304 32959
rect -6 32897 304 32931
rect -6 32869 42 32897
rect 70 32869 104 32897
rect 132 32869 166 32897
rect 194 32869 228 32897
rect 256 32869 304 32897
rect -6 32835 304 32869
rect -6 32807 42 32835
rect 70 32807 104 32835
rect 132 32807 166 32835
rect 194 32807 228 32835
rect 256 32807 304 32835
rect -6 32773 304 32807
rect -6 32745 42 32773
rect 70 32745 104 32773
rect 132 32745 166 32773
rect 194 32745 228 32773
rect 256 32745 304 32773
rect -6 23959 304 32745
rect -6 23931 42 23959
rect 70 23931 104 23959
rect 132 23931 166 23959
rect 194 23931 228 23959
rect 256 23931 304 23959
rect -6 23897 304 23931
rect -6 23869 42 23897
rect 70 23869 104 23897
rect 132 23869 166 23897
rect 194 23869 228 23897
rect 256 23869 304 23897
rect -6 23835 304 23869
rect -6 23807 42 23835
rect 70 23807 104 23835
rect 132 23807 166 23835
rect 194 23807 228 23835
rect 256 23807 304 23835
rect -6 23773 304 23807
rect -6 23745 42 23773
rect 70 23745 104 23773
rect 132 23745 166 23773
rect 194 23745 228 23773
rect 256 23745 304 23773
rect -6 14959 304 23745
rect -6 14931 42 14959
rect 70 14931 104 14959
rect 132 14931 166 14959
rect 194 14931 228 14959
rect 256 14931 304 14959
rect -6 14897 304 14931
rect -6 14869 42 14897
rect 70 14869 104 14897
rect 132 14869 166 14897
rect 194 14869 228 14897
rect 256 14869 304 14897
rect -6 14835 304 14869
rect -6 14807 42 14835
rect 70 14807 104 14835
rect 132 14807 166 14835
rect 194 14807 228 14835
rect 256 14807 304 14835
rect -6 14773 304 14807
rect -6 14745 42 14773
rect 70 14745 104 14773
rect 132 14745 166 14773
rect 194 14745 228 14773
rect 256 14745 304 14773
rect -6 5959 304 14745
rect -6 5931 42 5959
rect 70 5931 104 5959
rect 132 5931 166 5959
rect 194 5931 228 5959
rect 256 5931 304 5959
rect -6 5897 304 5931
rect -6 5869 42 5897
rect 70 5869 104 5897
rect 132 5869 166 5897
rect 194 5869 228 5897
rect 256 5869 304 5897
rect -6 5835 304 5869
rect -6 5807 42 5835
rect 70 5807 104 5835
rect 132 5807 166 5835
rect 194 5807 228 5835
rect 256 5807 304 5835
rect -6 5773 304 5807
rect -6 5745 42 5773
rect 70 5745 104 5773
rect 132 5745 166 5773
rect 194 5745 228 5773
rect 256 5745 304 5773
rect -6 424 304 5745
rect 474 299190 784 299238
rect 474 299162 522 299190
rect 550 299162 584 299190
rect 612 299162 646 299190
rect 674 299162 708 299190
rect 736 299162 784 299190
rect 474 299128 784 299162
rect 474 299100 522 299128
rect 550 299100 584 299128
rect 612 299100 646 299128
rect 674 299100 708 299128
rect 736 299100 784 299128
rect 474 299066 784 299100
rect 474 299038 522 299066
rect 550 299038 584 299066
rect 612 299038 646 299066
rect 674 299038 708 299066
rect 736 299038 784 299066
rect 474 299004 784 299038
rect 474 298976 522 299004
rect 550 298976 584 299004
rect 612 298976 646 299004
rect 674 298976 708 299004
rect 736 298976 784 299004
rect 474 290959 784 298976
rect 474 290931 522 290959
rect 550 290931 584 290959
rect 612 290931 646 290959
rect 674 290931 708 290959
rect 736 290931 784 290959
rect 474 290897 784 290931
rect 474 290869 522 290897
rect 550 290869 584 290897
rect 612 290869 646 290897
rect 674 290869 708 290897
rect 736 290869 784 290897
rect 474 290835 784 290869
rect 474 290807 522 290835
rect 550 290807 584 290835
rect 612 290807 646 290835
rect 674 290807 708 290835
rect 736 290807 784 290835
rect 474 290773 784 290807
rect 474 290745 522 290773
rect 550 290745 584 290773
rect 612 290745 646 290773
rect 674 290745 708 290773
rect 736 290745 784 290773
rect 474 281959 784 290745
rect 474 281931 522 281959
rect 550 281931 584 281959
rect 612 281931 646 281959
rect 674 281931 708 281959
rect 736 281931 784 281959
rect 474 281897 784 281931
rect 474 281869 522 281897
rect 550 281869 584 281897
rect 612 281869 646 281897
rect 674 281869 708 281897
rect 736 281869 784 281897
rect 474 281835 784 281869
rect 474 281807 522 281835
rect 550 281807 584 281835
rect 612 281807 646 281835
rect 674 281807 708 281835
rect 736 281807 784 281835
rect 474 281773 784 281807
rect 474 281745 522 281773
rect 550 281745 584 281773
rect 612 281745 646 281773
rect 674 281745 708 281773
rect 736 281745 784 281773
rect 474 272959 784 281745
rect 474 272931 522 272959
rect 550 272931 584 272959
rect 612 272931 646 272959
rect 674 272931 708 272959
rect 736 272931 784 272959
rect 474 272897 784 272931
rect 474 272869 522 272897
rect 550 272869 584 272897
rect 612 272869 646 272897
rect 674 272869 708 272897
rect 736 272869 784 272897
rect 474 272835 784 272869
rect 474 272807 522 272835
rect 550 272807 584 272835
rect 612 272807 646 272835
rect 674 272807 708 272835
rect 736 272807 784 272835
rect 474 272773 784 272807
rect 474 272745 522 272773
rect 550 272745 584 272773
rect 612 272745 646 272773
rect 674 272745 708 272773
rect 736 272745 784 272773
rect 474 263959 784 272745
rect 474 263931 522 263959
rect 550 263931 584 263959
rect 612 263931 646 263959
rect 674 263931 708 263959
rect 736 263931 784 263959
rect 474 263897 784 263931
rect 474 263869 522 263897
rect 550 263869 584 263897
rect 612 263869 646 263897
rect 674 263869 708 263897
rect 736 263869 784 263897
rect 474 263835 784 263869
rect 474 263807 522 263835
rect 550 263807 584 263835
rect 612 263807 646 263835
rect 674 263807 708 263835
rect 736 263807 784 263835
rect 474 263773 784 263807
rect 474 263745 522 263773
rect 550 263745 584 263773
rect 612 263745 646 263773
rect 674 263745 708 263773
rect 736 263745 784 263773
rect 474 254959 784 263745
rect 474 254931 522 254959
rect 550 254931 584 254959
rect 612 254931 646 254959
rect 674 254931 708 254959
rect 736 254931 784 254959
rect 474 254897 784 254931
rect 474 254869 522 254897
rect 550 254869 584 254897
rect 612 254869 646 254897
rect 674 254869 708 254897
rect 736 254869 784 254897
rect 474 254835 784 254869
rect 474 254807 522 254835
rect 550 254807 584 254835
rect 612 254807 646 254835
rect 674 254807 708 254835
rect 736 254807 784 254835
rect 474 254773 784 254807
rect 474 254745 522 254773
rect 550 254745 584 254773
rect 612 254745 646 254773
rect 674 254745 708 254773
rect 736 254745 784 254773
rect 474 245959 784 254745
rect 474 245931 522 245959
rect 550 245931 584 245959
rect 612 245931 646 245959
rect 674 245931 708 245959
rect 736 245931 784 245959
rect 474 245897 784 245931
rect 474 245869 522 245897
rect 550 245869 584 245897
rect 612 245869 646 245897
rect 674 245869 708 245897
rect 736 245869 784 245897
rect 474 245835 784 245869
rect 474 245807 522 245835
rect 550 245807 584 245835
rect 612 245807 646 245835
rect 674 245807 708 245835
rect 736 245807 784 245835
rect 474 245773 784 245807
rect 474 245745 522 245773
rect 550 245745 584 245773
rect 612 245745 646 245773
rect 674 245745 708 245773
rect 736 245745 784 245773
rect 474 236959 784 245745
rect 474 236931 522 236959
rect 550 236931 584 236959
rect 612 236931 646 236959
rect 674 236931 708 236959
rect 736 236931 784 236959
rect 474 236897 784 236931
rect 474 236869 522 236897
rect 550 236869 584 236897
rect 612 236869 646 236897
rect 674 236869 708 236897
rect 736 236869 784 236897
rect 474 236835 784 236869
rect 474 236807 522 236835
rect 550 236807 584 236835
rect 612 236807 646 236835
rect 674 236807 708 236835
rect 736 236807 784 236835
rect 474 236773 784 236807
rect 474 236745 522 236773
rect 550 236745 584 236773
rect 612 236745 646 236773
rect 674 236745 708 236773
rect 736 236745 784 236773
rect 474 227959 784 236745
rect 474 227931 522 227959
rect 550 227931 584 227959
rect 612 227931 646 227959
rect 674 227931 708 227959
rect 736 227931 784 227959
rect 474 227897 784 227931
rect 474 227869 522 227897
rect 550 227869 584 227897
rect 612 227869 646 227897
rect 674 227869 708 227897
rect 736 227869 784 227897
rect 474 227835 784 227869
rect 474 227807 522 227835
rect 550 227807 584 227835
rect 612 227807 646 227835
rect 674 227807 708 227835
rect 736 227807 784 227835
rect 474 227773 784 227807
rect 474 227745 522 227773
rect 550 227745 584 227773
rect 612 227745 646 227773
rect 674 227745 708 227773
rect 736 227745 784 227773
rect 474 218959 784 227745
rect 474 218931 522 218959
rect 550 218931 584 218959
rect 612 218931 646 218959
rect 674 218931 708 218959
rect 736 218931 784 218959
rect 474 218897 784 218931
rect 474 218869 522 218897
rect 550 218869 584 218897
rect 612 218869 646 218897
rect 674 218869 708 218897
rect 736 218869 784 218897
rect 474 218835 784 218869
rect 474 218807 522 218835
rect 550 218807 584 218835
rect 612 218807 646 218835
rect 674 218807 708 218835
rect 736 218807 784 218835
rect 474 218773 784 218807
rect 474 218745 522 218773
rect 550 218745 584 218773
rect 612 218745 646 218773
rect 674 218745 708 218773
rect 736 218745 784 218773
rect 474 209959 784 218745
rect 474 209931 522 209959
rect 550 209931 584 209959
rect 612 209931 646 209959
rect 674 209931 708 209959
rect 736 209931 784 209959
rect 474 209897 784 209931
rect 474 209869 522 209897
rect 550 209869 584 209897
rect 612 209869 646 209897
rect 674 209869 708 209897
rect 736 209869 784 209897
rect 474 209835 784 209869
rect 474 209807 522 209835
rect 550 209807 584 209835
rect 612 209807 646 209835
rect 674 209807 708 209835
rect 736 209807 784 209835
rect 474 209773 784 209807
rect 474 209745 522 209773
rect 550 209745 584 209773
rect 612 209745 646 209773
rect 674 209745 708 209773
rect 736 209745 784 209773
rect 474 200959 784 209745
rect 474 200931 522 200959
rect 550 200931 584 200959
rect 612 200931 646 200959
rect 674 200931 708 200959
rect 736 200931 784 200959
rect 474 200897 784 200931
rect 474 200869 522 200897
rect 550 200869 584 200897
rect 612 200869 646 200897
rect 674 200869 708 200897
rect 736 200869 784 200897
rect 474 200835 784 200869
rect 474 200807 522 200835
rect 550 200807 584 200835
rect 612 200807 646 200835
rect 674 200807 708 200835
rect 736 200807 784 200835
rect 474 200773 784 200807
rect 474 200745 522 200773
rect 550 200745 584 200773
rect 612 200745 646 200773
rect 674 200745 708 200773
rect 736 200745 784 200773
rect 474 191959 784 200745
rect 474 191931 522 191959
rect 550 191931 584 191959
rect 612 191931 646 191959
rect 674 191931 708 191959
rect 736 191931 784 191959
rect 474 191897 784 191931
rect 474 191869 522 191897
rect 550 191869 584 191897
rect 612 191869 646 191897
rect 674 191869 708 191897
rect 736 191869 784 191897
rect 474 191835 784 191869
rect 474 191807 522 191835
rect 550 191807 584 191835
rect 612 191807 646 191835
rect 674 191807 708 191835
rect 736 191807 784 191835
rect 474 191773 784 191807
rect 474 191745 522 191773
rect 550 191745 584 191773
rect 612 191745 646 191773
rect 674 191745 708 191773
rect 736 191745 784 191773
rect 474 182959 784 191745
rect 474 182931 522 182959
rect 550 182931 584 182959
rect 612 182931 646 182959
rect 674 182931 708 182959
rect 736 182931 784 182959
rect 474 182897 784 182931
rect 474 182869 522 182897
rect 550 182869 584 182897
rect 612 182869 646 182897
rect 674 182869 708 182897
rect 736 182869 784 182897
rect 474 182835 784 182869
rect 474 182807 522 182835
rect 550 182807 584 182835
rect 612 182807 646 182835
rect 674 182807 708 182835
rect 736 182807 784 182835
rect 474 182773 784 182807
rect 474 182745 522 182773
rect 550 182745 584 182773
rect 612 182745 646 182773
rect 674 182745 708 182773
rect 736 182745 784 182773
rect 474 173959 784 182745
rect 474 173931 522 173959
rect 550 173931 584 173959
rect 612 173931 646 173959
rect 674 173931 708 173959
rect 736 173931 784 173959
rect 474 173897 784 173931
rect 474 173869 522 173897
rect 550 173869 584 173897
rect 612 173869 646 173897
rect 674 173869 708 173897
rect 736 173869 784 173897
rect 474 173835 784 173869
rect 474 173807 522 173835
rect 550 173807 584 173835
rect 612 173807 646 173835
rect 674 173807 708 173835
rect 736 173807 784 173835
rect 474 173773 784 173807
rect 474 173745 522 173773
rect 550 173745 584 173773
rect 612 173745 646 173773
rect 674 173745 708 173773
rect 736 173745 784 173773
rect 474 164959 784 173745
rect 474 164931 522 164959
rect 550 164931 584 164959
rect 612 164931 646 164959
rect 674 164931 708 164959
rect 736 164931 784 164959
rect 474 164897 784 164931
rect 474 164869 522 164897
rect 550 164869 584 164897
rect 612 164869 646 164897
rect 674 164869 708 164897
rect 736 164869 784 164897
rect 474 164835 784 164869
rect 474 164807 522 164835
rect 550 164807 584 164835
rect 612 164807 646 164835
rect 674 164807 708 164835
rect 736 164807 784 164835
rect 474 164773 784 164807
rect 474 164745 522 164773
rect 550 164745 584 164773
rect 612 164745 646 164773
rect 674 164745 708 164773
rect 736 164745 784 164773
rect 474 155959 784 164745
rect 474 155931 522 155959
rect 550 155931 584 155959
rect 612 155931 646 155959
rect 674 155931 708 155959
rect 736 155931 784 155959
rect 474 155897 784 155931
rect 474 155869 522 155897
rect 550 155869 584 155897
rect 612 155869 646 155897
rect 674 155869 708 155897
rect 736 155869 784 155897
rect 474 155835 784 155869
rect 474 155807 522 155835
rect 550 155807 584 155835
rect 612 155807 646 155835
rect 674 155807 708 155835
rect 736 155807 784 155835
rect 474 155773 784 155807
rect 474 155745 522 155773
rect 550 155745 584 155773
rect 612 155745 646 155773
rect 674 155745 708 155773
rect 736 155745 784 155773
rect 474 146959 784 155745
rect 474 146931 522 146959
rect 550 146931 584 146959
rect 612 146931 646 146959
rect 674 146931 708 146959
rect 736 146931 784 146959
rect 474 146897 784 146931
rect 474 146869 522 146897
rect 550 146869 584 146897
rect 612 146869 646 146897
rect 674 146869 708 146897
rect 736 146869 784 146897
rect 474 146835 784 146869
rect 474 146807 522 146835
rect 550 146807 584 146835
rect 612 146807 646 146835
rect 674 146807 708 146835
rect 736 146807 784 146835
rect 474 146773 784 146807
rect 474 146745 522 146773
rect 550 146745 584 146773
rect 612 146745 646 146773
rect 674 146745 708 146773
rect 736 146745 784 146773
rect 474 137959 784 146745
rect 474 137931 522 137959
rect 550 137931 584 137959
rect 612 137931 646 137959
rect 674 137931 708 137959
rect 736 137931 784 137959
rect 474 137897 784 137931
rect 474 137869 522 137897
rect 550 137869 584 137897
rect 612 137869 646 137897
rect 674 137869 708 137897
rect 736 137869 784 137897
rect 474 137835 784 137869
rect 474 137807 522 137835
rect 550 137807 584 137835
rect 612 137807 646 137835
rect 674 137807 708 137835
rect 736 137807 784 137835
rect 474 137773 784 137807
rect 474 137745 522 137773
rect 550 137745 584 137773
rect 612 137745 646 137773
rect 674 137745 708 137773
rect 736 137745 784 137773
rect 474 128959 784 137745
rect 474 128931 522 128959
rect 550 128931 584 128959
rect 612 128931 646 128959
rect 674 128931 708 128959
rect 736 128931 784 128959
rect 474 128897 784 128931
rect 474 128869 522 128897
rect 550 128869 584 128897
rect 612 128869 646 128897
rect 674 128869 708 128897
rect 736 128869 784 128897
rect 474 128835 784 128869
rect 474 128807 522 128835
rect 550 128807 584 128835
rect 612 128807 646 128835
rect 674 128807 708 128835
rect 736 128807 784 128835
rect 474 128773 784 128807
rect 474 128745 522 128773
rect 550 128745 584 128773
rect 612 128745 646 128773
rect 674 128745 708 128773
rect 736 128745 784 128773
rect 474 119959 784 128745
rect 474 119931 522 119959
rect 550 119931 584 119959
rect 612 119931 646 119959
rect 674 119931 708 119959
rect 736 119931 784 119959
rect 474 119897 784 119931
rect 474 119869 522 119897
rect 550 119869 584 119897
rect 612 119869 646 119897
rect 674 119869 708 119897
rect 736 119869 784 119897
rect 474 119835 784 119869
rect 474 119807 522 119835
rect 550 119807 584 119835
rect 612 119807 646 119835
rect 674 119807 708 119835
rect 736 119807 784 119835
rect 474 119773 784 119807
rect 474 119745 522 119773
rect 550 119745 584 119773
rect 612 119745 646 119773
rect 674 119745 708 119773
rect 736 119745 784 119773
rect 474 110959 784 119745
rect 474 110931 522 110959
rect 550 110931 584 110959
rect 612 110931 646 110959
rect 674 110931 708 110959
rect 736 110931 784 110959
rect 474 110897 784 110931
rect 474 110869 522 110897
rect 550 110869 584 110897
rect 612 110869 646 110897
rect 674 110869 708 110897
rect 736 110869 784 110897
rect 474 110835 784 110869
rect 474 110807 522 110835
rect 550 110807 584 110835
rect 612 110807 646 110835
rect 674 110807 708 110835
rect 736 110807 784 110835
rect 474 110773 784 110807
rect 474 110745 522 110773
rect 550 110745 584 110773
rect 612 110745 646 110773
rect 674 110745 708 110773
rect 736 110745 784 110773
rect 474 101959 784 110745
rect 474 101931 522 101959
rect 550 101931 584 101959
rect 612 101931 646 101959
rect 674 101931 708 101959
rect 736 101931 784 101959
rect 474 101897 784 101931
rect 474 101869 522 101897
rect 550 101869 584 101897
rect 612 101869 646 101897
rect 674 101869 708 101897
rect 736 101869 784 101897
rect 474 101835 784 101869
rect 474 101807 522 101835
rect 550 101807 584 101835
rect 612 101807 646 101835
rect 674 101807 708 101835
rect 736 101807 784 101835
rect 474 101773 784 101807
rect 474 101745 522 101773
rect 550 101745 584 101773
rect 612 101745 646 101773
rect 674 101745 708 101773
rect 736 101745 784 101773
rect 474 92959 784 101745
rect 474 92931 522 92959
rect 550 92931 584 92959
rect 612 92931 646 92959
rect 674 92931 708 92959
rect 736 92931 784 92959
rect 474 92897 784 92931
rect 474 92869 522 92897
rect 550 92869 584 92897
rect 612 92869 646 92897
rect 674 92869 708 92897
rect 736 92869 784 92897
rect 474 92835 784 92869
rect 474 92807 522 92835
rect 550 92807 584 92835
rect 612 92807 646 92835
rect 674 92807 708 92835
rect 736 92807 784 92835
rect 474 92773 784 92807
rect 474 92745 522 92773
rect 550 92745 584 92773
rect 612 92745 646 92773
rect 674 92745 708 92773
rect 736 92745 784 92773
rect 474 83959 784 92745
rect 474 83931 522 83959
rect 550 83931 584 83959
rect 612 83931 646 83959
rect 674 83931 708 83959
rect 736 83931 784 83959
rect 474 83897 784 83931
rect 474 83869 522 83897
rect 550 83869 584 83897
rect 612 83869 646 83897
rect 674 83869 708 83897
rect 736 83869 784 83897
rect 474 83835 784 83869
rect 474 83807 522 83835
rect 550 83807 584 83835
rect 612 83807 646 83835
rect 674 83807 708 83835
rect 736 83807 784 83835
rect 474 83773 784 83807
rect 474 83745 522 83773
rect 550 83745 584 83773
rect 612 83745 646 83773
rect 674 83745 708 83773
rect 736 83745 784 83773
rect 474 74959 784 83745
rect 474 74931 522 74959
rect 550 74931 584 74959
rect 612 74931 646 74959
rect 674 74931 708 74959
rect 736 74931 784 74959
rect 474 74897 784 74931
rect 474 74869 522 74897
rect 550 74869 584 74897
rect 612 74869 646 74897
rect 674 74869 708 74897
rect 736 74869 784 74897
rect 474 74835 784 74869
rect 474 74807 522 74835
rect 550 74807 584 74835
rect 612 74807 646 74835
rect 674 74807 708 74835
rect 736 74807 784 74835
rect 474 74773 784 74807
rect 474 74745 522 74773
rect 550 74745 584 74773
rect 612 74745 646 74773
rect 674 74745 708 74773
rect 736 74745 784 74773
rect 474 65959 784 74745
rect 474 65931 522 65959
rect 550 65931 584 65959
rect 612 65931 646 65959
rect 674 65931 708 65959
rect 736 65931 784 65959
rect 474 65897 784 65931
rect 474 65869 522 65897
rect 550 65869 584 65897
rect 612 65869 646 65897
rect 674 65869 708 65897
rect 736 65869 784 65897
rect 474 65835 784 65869
rect 474 65807 522 65835
rect 550 65807 584 65835
rect 612 65807 646 65835
rect 674 65807 708 65835
rect 736 65807 784 65835
rect 474 65773 784 65807
rect 474 65745 522 65773
rect 550 65745 584 65773
rect 612 65745 646 65773
rect 674 65745 708 65773
rect 736 65745 784 65773
rect 474 56959 784 65745
rect 474 56931 522 56959
rect 550 56931 584 56959
rect 612 56931 646 56959
rect 674 56931 708 56959
rect 736 56931 784 56959
rect 474 56897 784 56931
rect 474 56869 522 56897
rect 550 56869 584 56897
rect 612 56869 646 56897
rect 674 56869 708 56897
rect 736 56869 784 56897
rect 474 56835 784 56869
rect 474 56807 522 56835
rect 550 56807 584 56835
rect 612 56807 646 56835
rect 674 56807 708 56835
rect 736 56807 784 56835
rect 474 56773 784 56807
rect 474 56745 522 56773
rect 550 56745 584 56773
rect 612 56745 646 56773
rect 674 56745 708 56773
rect 736 56745 784 56773
rect 474 47959 784 56745
rect 474 47931 522 47959
rect 550 47931 584 47959
rect 612 47931 646 47959
rect 674 47931 708 47959
rect 736 47931 784 47959
rect 474 47897 784 47931
rect 474 47869 522 47897
rect 550 47869 584 47897
rect 612 47869 646 47897
rect 674 47869 708 47897
rect 736 47869 784 47897
rect 474 47835 784 47869
rect 474 47807 522 47835
rect 550 47807 584 47835
rect 612 47807 646 47835
rect 674 47807 708 47835
rect 736 47807 784 47835
rect 474 47773 784 47807
rect 474 47745 522 47773
rect 550 47745 584 47773
rect 612 47745 646 47773
rect 674 47745 708 47773
rect 736 47745 784 47773
rect 474 38959 784 47745
rect 474 38931 522 38959
rect 550 38931 584 38959
rect 612 38931 646 38959
rect 674 38931 708 38959
rect 736 38931 784 38959
rect 474 38897 784 38931
rect 474 38869 522 38897
rect 550 38869 584 38897
rect 612 38869 646 38897
rect 674 38869 708 38897
rect 736 38869 784 38897
rect 474 38835 784 38869
rect 474 38807 522 38835
rect 550 38807 584 38835
rect 612 38807 646 38835
rect 674 38807 708 38835
rect 736 38807 784 38835
rect 474 38773 784 38807
rect 474 38745 522 38773
rect 550 38745 584 38773
rect 612 38745 646 38773
rect 674 38745 708 38773
rect 736 38745 784 38773
rect 474 29959 784 38745
rect 474 29931 522 29959
rect 550 29931 584 29959
rect 612 29931 646 29959
rect 674 29931 708 29959
rect 736 29931 784 29959
rect 474 29897 784 29931
rect 474 29869 522 29897
rect 550 29869 584 29897
rect 612 29869 646 29897
rect 674 29869 708 29897
rect 736 29869 784 29897
rect 474 29835 784 29869
rect 474 29807 522 29835
rect 550 29807 584 29835
rect 612 29807 646 29835
rect 674 29807 708 29835
rect 736 29807 784 29835
rect 474 29773 784 29807
rect 474 29745 522 29773
rect 550 29745 584 29773
rect 612 29745 646 29773
rect 674 29745 708 29773
rect 736 29745 784 29773
rect 474 20959 784 29745
rect 474 20931 522 20959
rect 550 20931 584 20959
rect 612 20931 646 20959
rect 674 20931 708 20959
rect 736 20931 784 20959
rect 474 20897 784 20931
rect 474 20869 522 20897
rect 550 20869 584 20897
rect 612 20869 646 20897
rect 674 20869 708 20897
rect 736 20869 784 20897
rect 474 20835 784 20869
rect 474 20807 522 20835
rect 550 20807 584 20835
rect 612 20807 646 20835
rect 674 20807 708 20835
rect 736 20807 784 20835
rect 474 20773 784 20807
rect 474 20745 522 20773
rect 550 20745 584 20773
rect 612 20745 646 20773
rect 674 20745 708 20773
rect 736 20745 784 20773
rect 474 11959 784 20745
rect 474 11931 522 11959
rect 550 11931 584 11959
rect 612 11931 646 11959
rect 674 11931 708 11959
rect 736 11931 784 11959
rect 474 11897 784 11931
rect 474 11869 522 11897
rect 550 11869 584 11897
rect 612 11869 646 11897
rect 674 11869 708 11897
rect 736 11869 784 11897
rect 474 11835 784 11869
rect 474 11807 522 11835
rect 550 11807 584 11835
rect 612 11807 646 11835
rect 674 11807 708 11835
rect 736 11807 784 11835
rect 474 11773 784 11807
rect 474 11745 522 11773
rect 550 11745 584 11773
rect 612 11745 646 11773
rect 674 11745 708 11773
rect 736 11745 784 11773
rect 474 2959 784 11745
rect 474 2931 522 2959
rect 550 2931 584 2959
rect 612 2931 646 2959
rect 674 2931 708 2959
rect 736 2931 784 2959
rect 474 2897 784 2931
rect 474 2869 522 2897
rect 550 2869 584 2897
rect 612 2869 646 2897
rect 674 2869 708 2897
rect 736 2869 784 2897
rect 474 2835 784 2869
rect 474 2807 522 2835
rect 550 2807 584 2835
rect 612 2807 646 2835
rect 674 2807 708 2835
rect 736 2807 784 2835
rect 474 2773 784 2807
rect 474 2745 522 2773
rect 550 2745 584 2773
rect 612 2745 646 2773
rect 674 2745 708 2773
rect 736 2745 784 2773
rect 474 904 784 2745
rect 474 876 522 904
rect 550 876 584 904
rect 612 876 646 904
rect 674 876 708 904
rect 736 876 784 904
rect 474 842 784 876
rect 474 814 522 842
rect 550 814 584 842
rect 612 814 646 842
rect 674 814 708 842
rect 736 814 784 842
rect 474 780 784 814
rect 474 752 522 780
rect 550 752 584 780
rect 612 752 646 780
rect 674 752 708 780
rect 736 752 784 780
rect 474 718 784 752
rect 474 690 522 718
rect 550 690 584 718
rect 612 690 646 718
rect 674 690 708 718
rect 736 690 784 718
rect 474 642 784 690
rect 2529 299190 2839 299718
rect 2529 299162 2577 299190
rect 2605 299162 2639 299190
rect 2667 299162 2701 299190
rect 2729 299162 2763 299190
rect 2791 299162 2839 299190
rect 2529 299128 2839 299162
rect 2529 299100 2577 299128
rect 2605 299100 2639 299128
rect 2667 299100 2701 299128
rect 2729 299100 2763 299128
rect 2791 299100 2839 299128
rect 2529 299066 2839 299100
rect 2529 299038 2577 299066
rect 2605 299038 2639 299066
rect 2667 299038 2701 299066
rect 2729 299038 2763 299066
rect 2791 299038 2839 299066
rect 2529 299004 2839 299038
rect 2529 298976 2577 299004
rect 2605 298976 2639 299004
rect 2667 298976 2701 299004
rect 2729 298976 2763 299004
rect 2791 298976 2839 299004
rect 2529 290959 2839 298976
rect 2529 290931 2577 290959
rect 2605 290931 2639 290959
rect 2667 290931 2701 290959
rect 2729 290931 2763 290959
rect 2791 290931 2839 290959
rect 2529 290897 2839 290931
rect 2529 290869 2577 290897
rect 2605 290869 2639 290897
rect 2667 290869 2701 290897
rect 2729 290869 2763 290897
rect 2791 290869 2839 290897
rect 2529 290835 2839 290869
rect 2529 290807 2577 290835
rect 2605 290807 2639 290835
rect 2667 290807 2701 290835
rect 2729 290807 2763 290835
rect 2791 290807 2839 290835
rect 2529 290773 2839 290807
rect 2529 290745 2577 290773
rect 2605 290745 2639 290773
rect 2667 290745 2701 290773
rect 2729 290745 2763 290773
rect 2791 290745 2839 290773
rect 2529 281959 2839 290745
rect 2529 281931 2577 281959
rect 2605 281931 2639 281959
rect 2667 281931 2701 281959
rect 2729 281931 2763 281959
rect 2791 281931 2839 281959
rect 2529 281897 2839 281931
rect 2529 281869 2577 281897
rect 2605 281869 2639 281897
rect 2667 281869 2701 281897
rect 2729 281869 2763 281897
rect 2791 281869 2839 281897
rect 2529 281835 2839 281869
rect 2529 281807 2577 281835
rect 2605 281807 2639 281835
rect 2667 281807 2701 281835
rect 2729 281807 2763 281835
rect 2791 281807 2839 281835
rect 2529 281773 2839 281807
rect 2529 281745 2577 281773
rect 2605 281745 2639 281773
rect 2667 281745 2701 281773
rect 2729 281745 2763 281773
rect 2791 281745 2839 281773
rect 2529 272959 2839 281745
rect 2529 272931 2577 272959
rect 2605 272931 2639 272959
rect 2667 272931 2701 272959
rect 2729 272931 2763 272959
rect 2791 272931 2839 272959
rect 2529 272897 2839 272931
rect 2529 272869 2577 272897
rect 2605 272869 2639 272897
rect 2667 272869 2701 272897
rect 2729 272869 2763 272897
rect 2791 272869 2839 272897
rect 2529 272835 2839 272869
rect 2529 272807 2577 272835
rect 2605 272807 2639 272835
rect 2667 272807 2701 272835
rect 2729 272807 2763 272835
rect 2791 272807 2839 272835
rect 2529 272773 2839 272807
rect 2529 272745 2577 272773
rect 2605 272745 2639 272773
rect 2667 272745 2701 272773
rect 2729 272745 2763 272773
rect 2791 272745 2839 272773
rect 2529 263959 2839 272745
rect 2529 263931 2577 263959
rect 2605 263931 2639 263959
rect 2667 263931 2701 263959
rect 2729 263931 2763 263959
rect 2791 263931 2839 263959
rect 2529 263897 2839 263931
rect 2529 263869 2577 263897
rect 2605 263869 2639 263897
rect 2667 263869 2701 263897
rect 2729 263869 2763 263897
rect 2791 263869 2839 263897
rect 2529 263835 2839 263869
rect 2529 263807 2577 263835
rect 2605 263807 2639 263835
rect 2667 263807 2701 263835
rect 2729 263807 2763 263835
rect 2791 263807 2839 263835
rect 2529 263773 2839 263807
rect 2529 263745 2577 263773
rect 2605 263745 2639 263773
rect 2667 263745 2701 263773
rect 2729 263745 2763 263773
rect 2791 263745 2839 263773
rect 2529 254959 2839 263745
rect 2529 254931 2577 254959
rect 2605 254931 2639 254959
rect 2667 254931 2701 254959
rect 2729 254931 2763 254959
rect 2791 254931 2839 254959
rect 2529 254897 2839 254931
rect 2529 254869 2577 254897
rect 2605 254869 2639 254897
rect 2667 254869 2701 254897
rect 2729 254869 2763 254897
rect 2791 254869 2839 254897
rect 2529 254835 2839 254869
rect 2529 254807 2577 254835
rect 2605 254807 2639 254835
rect 2667 254807 2701 254835
rect 2729 254807 2763 254835
rect 2791 254807 2839 254835
rect 2529 254773 2839 254807
rect 2529 254745 2577 254773
rect 2605 254745 2639 254773
rect 2667 254745 2701 254773
rect 2729 254745 2763 254773
rect 2791 254745 2839 254773
rect 2529 245959 2839 254745
rect 2529 245931 2577 245959
rect 2605 245931 2639 245959
rect 2667 245931 2701 245959
rect 2729 245931 2763 245959
rect 2791 245931 2839 245959
rect 2529 245897 2839 245931
rect 2529 245869 2577 245897
rect 2605 245869 2639 245897
rect 2667 245869 2701 245897
rect 2729 245869 2763 245897
rect 2791 245869 2839 245897
rect 2529 245835 2839 245869
rect 2529 245807 2577 245835
rect 2605 245807 2639 245835
rect 2667 245807 2701 245835
rect 2729 245807 2763 245835
rect 2791 245807 2839 245835
rect 2529 245773 2839 245807
rect 2529 245745 2577 245773
rect 2605 245745 2639 245773
rect 2667 245745 2701 245773
rect 2729 245745 2763 245773
rect 2791 245745 2839 245773
rect 2529 236959 2839 245745
rect 2529 236931 2577 236959
rect 2605 236931 2639 236959
rect 2667 236931 2701 236959
rect 2729 236931 2763 236959
rect 2791 236931 2839 236959
rect 2529 236897 2839 236931
rect 2529 236869 2577 236897
rect 2605 236869 2639 236897
rect 2667 236869 2701 236897
rect 2729 236869 2763 236897
rect 2791 236869 2839 236897
rect 2529 236835 2839 236869
rect 2529 236807 2577 236835
rect 2605 236807 2639 236835
rect 2667 236807 2701 236835
rect 2729 236807 2763 236835
rect 2791 236807 2839 236835
rect 2529 236773 2839 236807
rect 2529 236745 2577 236773
rect 2605 236745 2639 236773
rect 2667 236745 2701 236773
rect 2729 236745 2763 236773
rect 2791 236745 2839 236773
rect 2529 227959 2839 236745
rect 2529 227931 2577 227959
rect 2605 227931 2639 227959
rect 2667 227931 2701 227959
rect 2729 227931 2763 227959
rect 2791 227931 2839 227959
rect 2529 227897 2839 227931
rect 2529 227869 2577 227897
rect 2605 227869 2639 227897
rect 2667 227869 2701 227897
rect 2729 227869 2763 227897
rect 2791 227869 2839 227897
rect 2529 227835 2839 227869
rect 2529 227807 2577 227835
rect 2605 227807 2639 227835
rect 2667 227807 2701 227835
rect 2729 227807 2763 227835
rect 2791 227807 2839 227835
rect 2529 227773 2839 227807
rect 2529 227745 2577 227773
rect 2605 227745 2639 227773
rect 2667 227745 2701 227773
rect 2729 227745 2763 227773
rect 2791 227745 2839 227773
rect 2529 218959 2839 227745
rect 2529 218931 2577 218959
rect 2605 218931 2639 218959
rect 2667 218931 2701 218959
rect 2729 218931 2763 218959
rect 2791 218931 2839 218959
rect 2529 218897 2839 218931
rect 2529 218869 2577 218897
rect 2605 218869 2639 218897
rect 2667 218869 2701 218897
rect 2729 218869 2763 218897
rect 2791 218869 2839 218897
rect 2529 218835 2839 218869
rect 2529 218807 2577 218835
rect 2605 218807 2639 218835
rect 2667 218807 2701 218835
rect 2729 218807 2763 218835
rect 2791 218807 2839 218835
rect 2529 218773 2839 218807
rect 2529 218745 2577 218773
rect 2605 218745 2639 218773
rect 2667 218745 2701 218773
rect 2729 218745 2763 218773
rect 2791 218745 2839 218773
rect 2529 209959 2839 218745
rect 2529 209931 2577 209959
rect 2605 209931 2639 209959
rect 2667 209931 2701 209959
rect 2729 209931 2763 209959
rect 2791 209931 2839 209959
rect 2529 209897 2839 209931
rect 2529 209869 2577 209897
rect 2605 209869 2639 209897
rect 2667 209869 2701 209897
rect 2729 209869 2763 209897
rect 2791 209869 2839 209897
rect 2529 209835 2839 209869
rect 2529 209807 2577 209835
rect 2605 209807 2639 209835
rect 2667 209807 2701 209835
rect 2729 209807 2763 209835
rect 2791 209807 2839 209835
rect 2529 209773 2839 209807
rect 2529 209745 2577 209773
rect 2605 209745 2639 209773
rect 2667 209745 2701 209773
rect 2729 209745 2763 209773
rect 2791 209745 2839 209773
rect 2529 200959 2839 209745
rect 2529 200931 2577 200959
rect 2605 200931 2639 200959
rect 2667 200931 2701 200959
rect 2729 200931 2763 200959
rect 2791 200931 2839 200959
rect 2529 200897 2839 200931
rect 2529 200869 2577 200897
rect 2605 200869 2639 200897
rect 2667 200869 2701 200897
rect 2729 200869 2763 200897
rect 2791 200869 2839 200897
rect 2529 200835 2839 200869
rect 2529 200807 2577 200835
rect 2605 200807 2639 200835
rect 2667 200807 2701 200835
rect 2729 200807 2763 200835
rect 2791 200807 2839 200835
rect 2529 200773 2839 200807
rect 2529 200745 2577 200773
rect 2605 200745 2639 200773
rect 2667 200745 2701 200773
rect 2729 200745 2763 200773
rect 2791 200745 2839 200773
rect 2529 191959 2839 200745
rect 2529 191931 2577 191959
rect 2605 191931 2639 191959
rect 2667 191931 2701 191959
rect 2729 191931 2763 191959
rect 2791 191931 2839 191959
rect 2529 191897 2839 191931
rect 2529 191869 2577 191897
rect 2605 191869 2639 191897
rect 2667 191869 2701 191897
rect 2729 191869 2763 191897
rect 2791 191869 2839 191897
rect 2529 191835 2839 191869
rect 2529 191807 2577 191835
rect 2605 191807 2639 191835
rect 2667 191807 2701 191835
rect 2729 191807 2763 191835
rect 2791 191807 2839 191835
rect 2529 191773 2839 191807
rect 2529 191745 2577 191773
rect 2605 191745 2639 191773
rect 2667 191745 2701 191773
rect 2729 191745 2763 191773
rect 2791 191745 2839 191773
rect 2529 182959 2839 191745
rect 2529 182931 2577 182959
rect 2605 182931 2639 182959
rect 2667 182931 2701 182959
rect 2729 182931 2763 182959
rect 2791 182931 2839 182959
rect 2529 182897 2839 182931
rect 2529 182869 2577 182897
rect 2605 182869 2639 182897
rect 2667 182869 2701 182897
rect 2729 182869 2763 182897
rect 2791 182869 2839 182897
rect 2529 182835 2839 182869
rect 2529 182807 2577 182835
rect 2605 182807 2639 182835
rect 2667 182807 2701 182835
rect 2729 182807 2763 182835
rect 2791 182807 2839 182835
rect 2529 182773 2839 182807
rect 2529 182745 2577 182773
rect 2605 182745 2639 182773
rect 2667 182745 2701 182773
rect 2729 182745 2763 182773
rect 2791 182745 2839 182773
rect 2529 173959 2839 182745
rect 2529 173931 2577 173959
rect 2605 173931 2639 173959
rect 2667 173931 2701 173959
rect 2729 173931 2763 173959
rect 2791 173931 2839 173959
rect 2529 173897 2839 173931
rect 2529 173869 2577 173897
rect 2605 173869 2639 173897
rect 2667 173869 2701 173897
rect 2729 173869 2763 173897
rect 2791 173869 2839 173897
rect 2529 173835 2839 173869
rect 2529 173807 2577 173835
rect 2605 173807 2639 173835
rect 2667 173807 2701 173835
rect 2729 173807 2763 173835
rect 2791 173807 2839 173835
rect 2529 173773 2839 173807
rect 2529 173745 2577 173773
rect 2605 173745 2639 173773
rect 2667 173745 2701 173773
rect 2729 173745 2763 173773
rect 2791 173745 2839 173773
rect 2529 164959 2839 173745
rect 2529 164931 2577 164959
rect 2605 164931 2639 164959
rect 2667 164931 2701 164959
rect 2729 164931 2763 164959
rect 2791 164931 2839 164959
rect 2529 164897 2839 164931
rect 2529 164869 2577 164897
rect 2605 164869 2639 164897
rect 2667 164869 2701 164897
rect 2729 164869 2763 164897
rect 2791 164869 2839 164897
rect 2529 164835 2839 164869
rect 2529 164807 2577 164835
rect 2605 164807 2639 164835
rect 2667 164807 2701 164835
rect 2729 164807 2763 164835
rect 2791 164807 2839 164835
rect 2529 164773 2839 164807
rect 2529 164745 2577 164773
rect 2605 164745 2639 164773
rect 2667 164745 2701 164773
rect 2729 164745 2763 164773
rect 2791 164745 2839 164773
rect 2529 155959 2839 164745
rect 2529 155931 2577 155959
rect 2605 155931 2639 155959
rect 2667 155931 2701 155959
rect 2729 155931 2763 155959
rect 2791 155931 2839 155959
rect 2529 155897 2839 155931
rect 2529 155869 2577 155897
rect 2605 155869 2639 155897
rect 2667 155869 2701 155897
rect 2729 155869 2763 155897
rect 2791 155869 2839 155897
rect 2529 155835 2839 155869
rect 2529 155807 2577 155835
rect 2605 155807 2639 155835
rect 2667 155807 2701 155835
rect 2729 155807 2763 155835
rect 2791 155807 2839 155835
rect 2529 155773 2839 155807
rect 2529 155745 2577 155773
rect 2605 155745 2639 155773
rect 2667 155745 2701 155773
rect 2729 155745 2763 155773
rect 2791 155745 2839 155773
rect 2529 146959 2839 155745
rect 2529 146931 2577 146959
rect 2605 146931 2639 146959
rect 2667 146931 2701 146959
rect 2729 146931 2763 146959
rect 2791 146931 2839 146959
rect 2529 146897 2839 146931
rect 2529 146869 2577 146897
rect 2605 146869 2639 146897
rect 2667 146869 2701 146897
rect 2729 146869 2763 146897
rect 2791 146869 2839 146897
rect 2529 146835 2839 146869
rect 2529 146807 2577 146835
rect 2605 146807 2639 146835
rect 2667 146807 2701 146835
rect 2729 146807 2763 146835
rect 2791 146807 2839 146835
rect 2529 146773 2839 146807
rect 2529 146745 2577 146773
rect 2605 146745 2639 146773
rect 2667 146745 2701 146773
rect 2729 146745 2763 146773
rect 2791 146745 2839 146773
rect 2529 137959 2839 146745
rect 2529 137931 2577 137959
rect 2605 137931 2639 137959
rect 2667 137931 2701 137959
rect 2729 137931 2763 137959
rect 2791 137931 2839 137959
rect 2529 137897 2839 137931
rect 2529 137869 2577 137897
rect 2605 137869 2639 137897
rect 2667 137869 2701 137897
rect 2729 137869 2763 137897
rect 2791 137869 2839 137897
rect 2529 137835 2839 137869
rect 2529 137807 2577 137835
rect 2605 137807 2639 137835
rect 2667 137807 2701 137835
rect 2729 137807 2763 137835
rect 2791 137807 2839 137835
rect 2529 137773 2839 137807
rect 2529 137745 2577 137773
rect 2605 137745 2639 137773
rect 2667 137745 2701 137773
rect 2729 137745 2763 137773
rect 2791 137745 2839 137773
rect 2529 128959 2839 137745
rect 2529 128931 2577 128959
rect 2605 128931 2639 128959
rect 2667 128931 2701 128959
rect 2729 128931 2763 128959
rect 2791 128931 2839 128959
rect 2529 128897 2839 128931
rect 2529 128869 2577 128897
rect 2605 128869 2639 128897
rect 2667 128869 2701 128897
rect 2729 128869 2763 128897
rect 2791 128869 2839 128897
rect 2529 128835 2839 128869
rect 2529 128807 2577 128835
rect 2605 128807 2639 128835
rect 2667 128807 2701 128835
rect 2729 128807 2763 128835
rect 2791 128807 2839 128835
rect 2529 128773 2839 128807
rect 2529 128745 2577 128773
rect 2605 128745 2639 128773
rect 2667 128745 2701 128773
rect 2729 128745 2763 128773
rect 2791 128745 2839 128773
rect 2529 119959 2839 128745
rect 2529 119931 2577 119959
rect 2605 119931 2639 119959
rect 2667 119931 2701 119959
rect 2729 119931 2763 119959
rect 2791 119931 2839 119959
rect 2529 119897 2839 119931
rect 2529 119869 2577 119897
rect 2605 119869 2639 119897
rect 2667 119869 2701 119897
rect 2729 119869 2763 119897
rect 2791 119869 2839 119897
rect 2529 119835 2839 119869
rect 2529 119807 2577 119835
rect 2605 119807 2639 119835
rect 2667 119807 2701 119835
rect 2729 119807 2763 119835
rect 2791 119807 2839 119835
rect 2529 119773 2839 119807
rect 2529 119745 2577 119773
rect 2605 119745 2639 119773
rect 2667 119745 2701 119773
rect 2729 119745 2763 119773
rect 2791 119745 2839 119773
rect 2529 110959 2839 119745
rect 2529 110931 2577 110959
rect 2605 110931 2639 110959
rect 2667 110931 2701 110959
rect 2729 110931 2763 110959
rect 2791 110931 2839 110959
rect 2529 110897 2839 110931
rect 2529 110869 2577 110897
rect 2605 110869 2639 110897
rect 2667 110869 2701 110897
rect 2729 110869 2763 110897
rect 2791 110869 2839 110897
rect 2529 110835 2839 110869
rect 2529 110807 2577 110835
rect 2605 110807 2639 110835
rect 2667 110807 2701 110835
rect 2729 110807 2763 110835
rect 2791 110807 2839 110835
rect 2529 110773 2839 110807
rect 2529 110745 2577 110773
rect 2605 110745 2639 110773
rect 2667 110745 2701 110773
rect 2729 110745 2763 110773
rect 2791 110745 2839 110773
rect 2529 101959 2839 110745
rect 2529 101931 2577 101959
rect 2605 101931 2639 101959
rect 2667 101931 2701 101959
rect 2729 101931 2763 101959
rect 2791 101931 2839 101959
rect 2529 101897 2839 101931
rect 2529 101869 2577 101897
rect 2605 101869 2639 101897
rect 2667 101869 2701 101897
rect 2729 101869 2763 101897
rect 2791 101869 2839 101897
rect 2529 101835 2839 101869
rect 2529 101807 2577 101835
rect 2605 101807 2639 101835
rect 2667 101807 2701 101835
rect 2729 101807 2763 101835
rect 2791 101807 2839 101835
rect 2529 101773 2839 101807
rect 2529 101745 2577 101773
rect 2605 101745 2639 101773
rect 2667 101745 2701 101773
rect 2729 101745 2763 101773
rect 2791 101745 2839 101773
rect 2529 92959 2839 101745
rect 2529 92931 2577 92959
rect 2605 92931 2639 92959
rect 2667 92931 2701 92959
rect 2729 92931 2763 92959
rect 2791 92931 2839 92959
rect 2529 92897 2839 92931
rect 2529 92869 2577 92897
rect 2605 92869 2639 92897
rect 2667 92869 2701 92897
rect 2729 92869 2763 92897
rect 2791 92869 2839 92897
rect 2529 92835 2839 92869
rect 2529 92807 2577 92835
rect 2605 92807 2639 92835
rect 2667 92807 2701 92835
rect 2729 92807 2763 92835
rect 2791 92807 2839 92835
rect 2529 92773 2839 92807
rect 2529 92745 2577 92773
rect 2605 92745 2639 92773
rect 2667 92745 2701 92773
rect 2729 92745 2763 92773
rect 2791 92745 2839 92773
rect 2529 83959 2839 92745
rect 2529 83931 2577 83959
rect 2605 83931 2639 83959
rect 2667 83931 2701 83959
rect 2729 83931 2763 83959
rect 2791 83931 2839 83959
rect 2529 83897 2839 83931
rect 2529 83869 2577 83897
rect 2605 83869 2639 83897
rect 2667 83869 2701 83897
rect 2729 83869 2763 83897
rect 2791 83869 2839 83897
rect 2529 83835 2839 83869
rect 2529 83807 2577 83835
rect 2605 83807 2639 83835
rect 2667 83807 2701 83835
rect 2729 83807 2763 83835
rect 2791 83807 2839 83835
rect 2529 83773 2839 83807
rect 2529 83745 2577 83773
rect 2605 83745 2639 83773
rect 2667 83745 2701 83773
rect 2729 83745 2763 83773
rect 2791 83745 2839 83773
rect 2529 74959 2839 83745
rect 2529 74931 2577 74959
rect 2605 74931 2639 74959
rect 2667 74931 2701 74959
rect 2729 74931 2763 74959
rect 2791 74931 2839 74959
rect 2529 74897 2839 74931
rect 2529 74869 2577 74897
rect 2605 74869 2639 74897
rect 2667 74869 2701 74897
rect 2729 74869 2763 74897
rect 2791 74869 2839 74897
rect 2529 74835 2839 74869
rect 2529 74807 2577 74835
rect 2605 74807 2639 74835
rect 2667 74807 2701 74835
rect 2729 74807 2763 74835
rect 2791 74807 2839 74835
rect 2529 74773 2839 74807
rect 2529 74745 2577 74773
rect 2605 74745 2639 74773
rect 2667 74745 2701 74773
rect 2729 74745 2763 74773
rect 2791 74745 2839 74773
rect 2529 65959 2839 74745
rect 2529 65931 2577 65959
rect 2605 65931 2639 65959
rect 2667 65931 2701 65959
rect 2729 65931 2763 65959
rect 2791 65931 2839 65959
rect 2529 65897 2839 65931
rect 2529 65869 2577 65897
rect 2605 65869 2639 65897
rect 2667 65869 2701 65897
rect 2729 65869 2763 65897
rect 2791 65869 2839 65897
rect 2529 65835 2839 65869
rect 2529 65807 2577 65835
rect 2605 65807 2639 65835
rect 2667 65807 2701 65835
rect 2729 65807 2763 65835
rect 2791 65807 2839 65835
rect 2529 65773 2839 65807
rect 2529 65745 2577 65773
rect 2605 65745 2639 65773
rect 2667 65745 2701 65773
rect 2729 65745 2763 65773
rect 2791 65745 2839 65773
rect 2529 56959 2839 65745
rect 2529 56931 2577 56959
rect 2605 56931 2639 56959
rect 2667 56931 2701 56959
rect 2729 56931 2763 56959
rect 2791 56931 2839 56959
rect 2529 56897 2839 56931
rect 2529 56869 2577 56897
rect 2605 56869 2639 56897
rect 2667 56869 2701 56897
rect 2729 56869 2763 56897
rect 2791 56869 2839 56897
rect 2529 56835 2839 56869
rect 2529 56807 2577 56835
rect 2605 56807 2639 56835
rect 2667 56807 2701 56835
rect 2729 56807 2763 56835
rect 2791 56807 2839 56835
rect 2529 56773 2839 56807
rect 2529 56745 2577 56773
rect 2605 56745 2639 56773
rect 2667 56745 2701 56773
rect 2729 56745 2763 56773
rect 2791 56745 2839 56773
rect 2529 47959 2839 56745
rect 2529 47931 2577 47959
rect 2605 47931 2639 47959
rect 2667 47931 2701 47959
rect 2729 47931 2763 47959
rect 2791 47931 2839 47959
rect 2529 47897 2839 47931
rect 2529 47869 2577 47897
rect 2605 47869 2639 47897
rect 2667 47869 2701 47897
rect 2729 47869 2763 47897
rect 2791 47869 2839 47897
rect 2529 47835 2839 47869
rect 2529 47807 2577 47835
rect 2605 47807 2639 47835
rect 2667 47807 2701 47835
rect 2729 47807 2763 47835
rect 2791 47807 2839 47835
rect 2529 47773 2839 47807
rect 2529 47745 2577 47773
rect 2605 47745 2639 47773
rect 2667 47745 2701 47773
rect 2729 47745 2763 47773
rect 2791 47745 2839 47773
rect 2529 38959 2839 47745
rect 2529 38931 2577 38959
rect 2605 38931 2639 38959
rect 2667 38931 2701 38959
rect 2729 38931 2763 38959
rect 2791 38931 2839 38959
rect 2529 38897 2839 38931
rect 2529 38869 2577 38897
rect 2605 38869 2639 38897
rect 2667 38869 2701 38897
rect 2729 38869 2763 38897
rect 2791 38869 2839 38897
rect 2529 38835 2839 38869
rect 2529 38807 2577 38835
rect 2605 38807 2639 38835
rect 2667 38807 2701 38835
rect 2729 38807 2763 38835
rect 2791 38807 2839 38835
rect 2529 38773 2839 38807
rect 2529 38745 2577 38773
rect 2605 38745 2639 38773
rect 2667 38745 2701 38773
rect 2729 38745 2763 38773
rect 2791 38745 2839 38773
rect 2529 29959 2839 38745
rect 2529 29931 2577 29959
rect 2605 29931 2639 29959
rect 2667 29931 2701 29959
rect 2729 29931 2763 29959
rect 2791 29931 2839 29959
rect 2529 29897 2839 29931
rect 2529 29869 2577 29897
rect 2605 29869 2639 29897
rect 2667 29869 2701 29897
rect 2729 29869 2763 29897
rect 2791 29869 2839 29897
rect 2529 29835 2839 29869
rect 2529 29807 2577 29835
rect 2605 29807 2639 29835
rect 2667 29807 2701 29835
rect 2729 29807 2763 29835
rect 2791 29807 2839 29835
rect 2529 29773 2839 29807
rect 2529 29745 2577 29773
rect 2605 29745 2639 29773
rect 2667 29745 2701 29773
rect 2729 29745 2763 29773
rect 2791 29745 2839 29773
rect 2529 20959 2839 29745
rect 2529 20931 2577 20959
rect 2605 20931 2639 20959
rect 2667 20931 2701 20959
rect 2729 20931 2763 20959
rect 2791 20931 2839 20959
rect 2529 20897 2839 20931
rect 2529 20869 2577 20897
rect 2605 20869 2639 20897
rect 2667 20869 2701 20897
rect 2729 20869 2763 20897
rect 2791 20869 2839 20897
rect 2529 20835 2839 20869
rect 2529 20807 2577 20835
rect 2605 20807 2639 20835
rect 2667 20807 2701 20835
rect 2729 20807 2763 20835
rect 2791 20807 2839 20835
rect 2529 20773 2839 20807
rect 2529 20745 2577 20773
rect 2605 20745 2639 20773
rect 2667 20745 2701 20773
rect 2729 20745 2763 20773
rect 2791 20745 2839 20773
rect 2529 11959 2839 20745
rect 2529 11931 2577 11959
rect 2605 11931 2639 11959
rect 2667 11931 2701 11959
rect 2729 11931 2763 11959
rect 2791 11931 2839 11959
rect 2529 11897 2839 11931
rect 2529 11869 2577 11897
rect 2605 11869 2639 11897
rect 2667 11869 2701 11897
rect 2729 11869 2763 11897
rect 2791 11869 2839 11897
rect 2529 11835 2839 11869
rect 2529 11807 2577 11835
rect 2605 11807 2639 11835
rect 2667 11807 2701 11835
rect 2729 11807 2763 11835
rect 2791 11807 2839 11835
rect 2529 11773 2839 11807
rect 2529 11745 2577 11773
rect 2605 11745 2639 11773
rect 2667 11745 2701 11773
rect 2729 11745 2763 11773
rect 2791 11745 2839 11773
rect 2529 2959 2839 11745
rect 2529 2931 2577 2959
rect 2605 2931 2639 2959
rect 2667 2931 2701 2959
rect 2729 2931 2763 2959
rect 2791 2931 2839 2959
rect 2529 2897 2839 2931
rect 2529 2869 2577 2897
rect 2605 2869 2639 2897
rect 2667 2869 2701 2897
rect 2729 2869 2763 2897
rect 2791 2869 2839 2897
rect 2529 2835 2839 2869
rect 2529 2807 2577 2835
rect 2605 2807 2639 2835
rect 2667 2807 2701 2835
rect 2729 2807 2763 2835
rect 2791 2807 2839 2835
rect 2529 2773 2839 2807
rect 2529 2745 2577 2773
rect 2605 2745 2639 2773
rect 2667 2745 2701 2773
rect 2729 2745 2763 2773
rect 2791 2745 2839 2773
rect 2529 904 2839 2745
rect 2529 876 2577 904
rect 2605 876 2639 904
rect 2667 876 2701 904
rect 2729 876 2763 904
rect 2791 876 2839 904
rect 2529 842 2839 876
rect 2529 814 2577 842
rect 2605 814 2639 842
rect 2667 814 2701 842
rect 2729 814 2763 842
rect 2791 814 2839 842
rect 2529 780 2839 814
rect 2529 752 2577 780
rect 2605 752 2639 780
rect 2667 752 2701 780
rect 2729 752 2763 780
rect 2791 752 2839 780
rect 2529 718 2839 752
rect 2529 690 2577 718
rect 2605 690 2639 718
rect 2667 690 2701 718
rect 2729 690 2763 718
rect 2791 690 2839 718
rect -6 396 42 424
rect 70 396 104 424
rect 132 396 166 424
rect 194 396 228 424
rect 256 396 304 424
rect -6 362 304 396
rect -6 334 42 362
rect 70 334 104 362
rect 132 334 166 362
rect 194 334 228 362
rect 256 334 304 362
rect -6 300 304 334
rect -6 272 42 300
rect 70 272 104 300
rect 132 272 166 300
rect 194 272 228 300
rect 256 272 304 300
rect -6 238 304 272
rect -6 210 42 238
rect 70 210 104 238
rect 132 210 166 238
rect 194 210 228 238
rect 256 210 304 238
rect -6 162 304 210
rect 2529 162 2839 690
rect 4389 299670 4699 299718
rect 4389 299642 4437 299670
rect 4465 299642 4499 299670
rect 4527 299642 4561 299670
rect 4589 299642 4623 299670
rect 4651 299642 4699 299670
rect 4389 299608 4699 299642
rect 4389 299580 4437 299608
rect 4465 299580 4499 299608
rect 4527 299580 4561 299608
rect 4589 299580 4623 299608
rect 4651 299580 4699 299608
rect 4389 299546 4699 299580
rect 4389 299518 4437 299546
rect 4465 299518 4499 299546
rect 4527 299518 4561 299546
rect 4589 299518 4623 299546
rect 4651 299518 4699 299546
rect 4389 299484 4699 299518
rect 4389 299456 4437 299484
rect 4465 299456 4499 299484
rect 4527 299456 4561 299484
rect 4589 299456 4623 299484
rect 4651 299456 4699 299484
rect 4389 293959 4699 299456
rect 4389 293931 4437 293959
rect 4465 293931 4499 293959
rect 4527 293931 4561 293959
rect 4589 293931 4623 293959
rect 4651 293931 4699 293959
rect 4389 293897 4699 293931
rect 4389 293869 4437 293897
rect 4465 293869 4499 293897
rect 4527 293869 4561 293897
rect 4589 293869 4623 293897
rect 4651 293869 4699 293897
rect 4389 293835 4699 293869
rect 4389 293807 4437 293835
rect 4465 293807 4499 293835
rect 4527 293807 4561 293835
rect 4589 293807 4623 293835
rect 4651 293807 4699 293835
rect 4389 293773 4699 293807
rect 4389 293745 4437 293773
rect 4465 293745 4499 293773
rect 4527 293745 4561 293773
rect 4589 293745 4623 293773
rect 4651 293745 4699 293773
rect 4389 284959 4699 293745
rect 4389 284931 4437 284959
rect 4465 284931 4499 284959
rect 4527 284931 4561 284959
rect 4589 284931 4623 284959
rect 4651 284931 4699 284959
rect 4389 284897 4699 284931
rect 4389 284869 4437 284897
rect 4465 284869 4499 284897
rect 4527 284869 4561 284897
rect 4589 284869 4623 284897
rect 4651 284869 4699 284897
rect 4389 284835 4699 284869
rect 4389 284807 4437 284835
rect 4465 284807 4499 284835
rect 4527 284807 4561 284835
rect 4589 284807 4623 284835
rect 4651 284807 4699 284835
rect 4389 284773 4699 284807
rect 4389 284745 4437 284773
rect 4465 284745 4499 284773
rect 4527 284745 4561 284773
rect 4589 284745 4623 284773
rect 4651 284745 4699 284773
rect 4389 275959 4699 284745
rect 4389 275931 4437 275959
rect 4465 275931 4499 275959
rect 4527 275931 4561 275959
rect 4589 275931 4623 275959
rect 4651 275931 4699 275959
rect 4389 275897 4699 275931
rect 4389 275869 4437 275897
rect 4465 275869 4499 275897
rect 4527 275869 4561 275897
rect 4589 275869 4623 275897
rect 4651 275869 4699 275897
rect 4389 275835 4699 275869
rect 4389 275807 4437 275835
rect 4465 275807 4499 275835
rect 4527 275807 4561 275835
rect 4589 275807 4623 275835
rect 4651 275807 4699 275835
rect 4389 275773 4699 275807
rect 4389 275745 4437 275773
rect 4465 275745 4499 275773
rect 4527 275745 4561 275773
rect 4589 275745 4623 275773
rect 4651 275745 4699 275773
rect 4389 266959 4699 275745
rect 4389 266931 4437 266959
rect 4465 266931 4499 266959
rect 4527 266931 4561 266959
rect 4589 266931 4623 266959
rect 4651 266931 4699 266959
rect 4389 266897 4699 266931
rect 4389 266869 4437 266897
rect 4465 266869 4499 266897
rect 4527 266869 4561 266897
rect 4589 266869 4623 266897
rect 4651 266869 4699 266897
rect 4389 266835 4699 266869
rect 4389 266807 4437 266835
rect 4465 266807 4499 266835
rect 4527 266807 4561 266835
rect 4589 266807 4623 266835
rect 4651 266807 4699 266835
rect 4389 266773 4699 266807
rect 4389 266745 4437 266773
rect 4465 266745 4499 266773
rect 4527 266745 4561 266773
rect 4589 266745 4623 266773
rect 4651 266745 4699 266773
rect 4389 257959 4699 266745
rect 4389 257931 4437 257959
rect 4465 257931 4499 257959
rect 4527 257931 4561 257959
rect 4589 257931 4623 257959
rect 4651 257931 4699 257959
rect 4389 257897 4699 257931
rect 4389 257869 4437 257897
rect 4465 257869 4499 257897
rect 4527 257869 4561 257897
rect 4589 257869 4623 257897
rect 4651 257869 4699 257897
rect 4389 257835 4699 257869
rect 4389 257807 4437 257835
rect 4465 257807 4499 257835
rect 4527 257807 4561 257835
rect 4589 257807 4623 257835
rect 4651 257807 4699 257835
rect 4389 257773 4699 257807
rect 4389 257745 4437 257773
rect 4465 257745 4499 257773
rect 4527 257745 4561 257773
rect 4589 257745 4623 257773
rect 4651 257745 4699 257773
rect 4389 248959 4699 257745
rect 4389 248931 4437 248959
rect 4465 248931 4499 248959
rect 4527 248931 4561 248959
rect 4589 248931 4623 248959
rect 4651 248931 4699 248959
rect 4389 248897 4699 248931
rect 4389 248869 4437 248897
rect 4465 248869 4499 248897
rect 4527 248869 4561 248897
rect 4589 248869 4623 248897
rect 4651 248869 4699 248897
rect 4389 248835 4699 248869
rect 4389 248807 4437 248835
rect 4465 248807 4499 248835
rect 4527 248807 4561 248835
rect 4589 248807 4623 248835
rect 4651 248807 4699 248835
rect 4389 248773 4699 248807
rect 4389 248745 4437 248773
rect 4465 248745 4499 248773
rect 4527 248745 4561 248773
rect 4589 248745 4623 248773
rect 4651 248745 4699 248773
rect 4389 239959 4699 248745
rect 4389 239931 4437 239959
rect 4465 239931 4499 239959
rect 4527 239931 4561 239959
rect 4589 239931 4623 239959
rect 4651 239931 4699 239959
rect 4389 239897 4699 239931
rect 4389 239869 4437 239897
rect 4465 239869 4499 239897
rect 4527 239869 4561 239897
rect 4589 239869 4623 239897
rect 4651 239869 4699 239897
rect 4389 239835 4699 239869
rect 4389 239807 4437 239835
rect 4465 239807 4499 239835
rect 4527 239807 4561 239835
rect 4589 239807 4623 239835
rect 4651 239807 4699 239835
rect 4389 239773 4699 239807
rect 4389 239745 4437 239773
rect 4465 239745 4499 239773
rect 4527 239745 4561 239773
rect 4589 239745 4623 239773
rect 4651 239745 4699 239773
rect 4389 230959 4699 239745
rect 4389 230931 4437 230959
rect 4465 230931 4499 230959
rect 4527 230931 4561 230959
rect 4589 230931 4623 230959
rect 4651 230931 4699 230959
rect 4389 230897 4699 230931
rect 4389 230869 4437 230897
rect 4465 230869 4499 230897
rect 4527 230869 4561 230897
rect 4589 230869 4623 230897
rect 4651 230869 4699 230897
rect 4389 230835 4699 230869
rect 4389 230807 4437 230835
rect 4465 230807 4499 230835
rect 4527 230807 4561 230835
rect 4589 230807 4623 230835
rect 4651 230807 4699 230835
rect 4389 230773 4699 230807
rect 4389 230745 4437 230773
rect 4465 230745 4499 230773
rect 4527 230745 4561 230773
rect 4589 230745 4623 230773
rect 4651 230745 4699 230773
rect 4389 221959 4699 230745
rect 4389 221931 4437 221959
rect 4465 221931 4499 221959
rect 4527 221931 4561 221959
rect 4589 221931 4623 221959
rect 4651 221931 4699 221959
rect 4389 221897 4699 221931
rect 4389 221869 4437 221897
rect 4465 221869 4499 221897
rect 4527 221869 4561 221897
rect 4589 221869 4623 221897
rect 4651 221869 4699 221897
rect 4389 221835 4699 221869
rect 4389 221807 4437 221835
rect 4465 221807 4499 221835
rect 4527 221807 4561 221835
rect 4589 221807 4623 221835
rect 4651 221807 4699 221835
rect 4389 221773 4699 221807
rect 4389 221745 4437 221773
rect 4465 221745 4499 221773
rect 4527 221745 4561 221773
rect 4589 221745 4623 221773
rect 4651 221745 4699 221773
rect 4389 212959 4699 221745
rect 4389 212931 4437 212959
rect 4465 212931 4499 212959
rect 4527 212931 4561 212959
rect 4589 212931 4623 212959
rect 4651 212931 4699 212959
rect 4389 212897 4699 212931
rect 4389 212869 4437 212897
rect 4465 212869 4499 212897
rect 4527 212869 4561 212897
rect 4589 212869 4623 212897
rect 4651 212869 4699 212897
rect 4389 212835 4699 212869
rect 4389 212807 4437 212835
rect 4465 212807 4499 212835
rect 4527 212807 4561 212835
rect 4589 212807 4623 212835
rect 4651 212807 4699 212835
rect 4389 212773 4699 212807
rect 4389 212745 4437 212773
rect 4465 212745 4499 212773
rect 4527 212745 4561 212773
rect 4589 212745 4623 212773
rect 4651 212745 4699 212773
rect 4389 203959 4699 212745
rect 4389 203931 4437 203959
rect 4465 203931 4499 203959
rect 4527 203931 4561 203959
rect 4589 203931 4623 203959
rect 4651 203931 4699 203959
rect 4389 203897 4699 203931
rect 4389 203869 4437 203897
rect 4465 203869 4499 203897
rect 4527 203869 4561 203897
rect 4589 203869 4623 203897
rect 4651 203869 4699 203897
rect 4389 203835 4699 203869
rect 4389 203807 4437 203835
rect 4465 203807 4499 203835
rect 4527 203807 4561 203835
rect 4589 203807 4623 203835
rect 4651 203807 4699 203835
rect 4389 203773 4699 203807
rect 4389 203745 4437 203773
rect 4465 203745 4499 203773
rect 4527 203745 4561 203773
rect 4589 203745 4623 203773
rect 4651 203745 4699 203773
rect 4389 194959 4699 203745
rect 4389 194931 4437 194959
rect 4465 194931 4499 194959
rect 4527 194931 4561 194959
rect 4589 194931 4623 194959
rect 4651 194931 4699 194959
rect 4389 194897 4699 194931
rect 4389 194869 4437 194897
rect 4465 194869 4499 194897
rect 4527 194869 4561 194897
rect 4589 194869 4623 194897
rect 4651 194869 4699 194897
rect 4389 194835 4699 194869
rect 4389 194807 4437 194835
rect 4465 194807 4499 194835
rect 4527 194807 4561 194835
rect 4589 194807 4623 194835
rect 4651 194807 4699 194835
rect 4389 194773 4699 194807
rect 4389 194745 4437 194773
rect 4465 194745 4499 194773
rect 4527 194745 4561 194773
rect 4589 194745 4623 194773
rect 4651 194745 4699 194773
rect 4389 185959 4699 194745
rect 4389 185931 4437 185959
rect 4465 185931 4499 185959
rect 4527 185931 4561 185959
rect 4589 185931 4623 185959
rect 4651 185931 4699 185959
rect 4389 185897 4699 185931
rect 4389 185869 4437 185897
rect 4465 185869 4499 185897
rect 4527 185869 4561 185897
rect 4589 185869 4623 185897
rect 4651 185869 4699 185897
rect 4389 185835 4699 185869
rect 4389 185807 4437 185835
rect 4465 185807 4499 185835
rect 4527 185807 4561 185835
rect 4589 185807 4623 185835
rect 4651 185807 4699 185835
rect 4389 185773 4699 185807
rect 4389 185745 4437 185773
rect 4465 185745 4499 185773
rect 4527 185745 4561 185773
rect 4589 185745 4623 185773
rect 4651 185745 4699 185773
rect 4389 176959 4699 185745
rect 4389 176931 4437 176959
rect 4465 176931 4499 176959
rect 4527 176931 4561 176959
rect 4589 176931 4623 176959
rect 4651 176931 4699 176959
rect 4389 176897 4699 176931
rect 4389 176869 4437 176897
rect 4465 176869 4499 176897
rect 4527 176869 4561 176897
rect 4589 176869 4623 176897
rect 4651 176869 4699 176897
rect 4389 176835 4699 176869
rect 4389 176807 4437 176835
rect 4465 176807 4499 176835
rect 4527 176807 4561 176835
rect 4589 176807 4623 176835
rect 4651 176807 4699 176835
rect 4389 176773 4699 176807
rect 4389 176745 4437 176773
rect 4465 176745 4499 176773
rect 4527 176745 4561 176773
rect 4589 176745 4623 176773
rect 4651 176745 4699 176773
rect 4389 167959 4699 176745
rect 4389 167931 4437 167959
rect 4465 167931 4499 167959
rect 4527 167931 4561 167959
rect 4589 167931 4623 167959
rect 4651 167931 4699 167959
rect 4389 167897 4699 167931
rect 4389 167869 4437 167897
rect 4465 167869 4499 167897
rect 4527 167869 4561 167897
rect 4589 167869 4623 167897
rect 4651 167869 4699 167897
rect 4389 167835 4699 167869
rect 4389 167807 4437 167835
rect 4465 167807 4499 167835
rect 4527 167807 4561 167835
rect 4589 167807 4623 167835
rect 4651 167807 4699 167835
rect 4389 167773 4699 167807
rect 4389 167745 4437 167773
rect 4465 167745 4499 167773
rect 4527 167745 4561 167773
rect 4589 167745 4623 167773
rect 4651 167745 4699 167773
rect 4389 158959 4699 167745
rect 4389 158931 4437 158959
rect 4465 158931 4499 158959
rect 4527 158931 4561 158959
rect 4589 158931 4623 158959
rect 4651 158931 4699 158959
rect 4389 158897 4699 158931
rect 4389 158869 4437 158897
rect 4465 158869 4499 158897
rect 4527 158869 4561 158897
rect 4589 158869 4623 158897
rect 4651 158869 4699 158897
rect 4389 158835 4699 158869
rect 4389 158807 4437 158835
rect 4465 158807 4499 158835
rect 4527 158807 4561 158835
rect 4589 158807 4623 158835
rect 4651 158807 4699 158835
rect 4389 158773 4699 158807
rect 4389 158745 4437 158773
rect 4465 158745 4499 158773
rect 4527 158745 4561 158773
rect 4589 158745 4623 158773
rect 4651 158745 4699 158773
rect 4389 149959 4699 158745
rect 4389 149931 4437 149959
rect 4465 149931 4499 149959
rect 4527 149931 4561 149959
rect 4589 149931 4623 149959
rect 4651 149931 4699 149959
rect 4389 149897 4699 149931
rect 4389 149869 4437 149897
rect 4465 149869 4499 149897
rect 4527 149869 4561 149897
rect 4589 149869 4623 149897
rect 4651 149869 4699 149897
rect 4389 149835 4699 149869
rect 4389 149807 4437 149835
rect 4465 149807 4499 149835
rect 4527 149807 4561 149835
rect 4589 149807 4623 149835
rect 4651 149807 4699 149835
rect 4389 149773 4699 149807
rect 4389 149745 4437 149773
rect 4465 149745 4499 149773
rect 4527 149745 4561 149773
rect 4589 149745 4623 149773
rect 4651 149745 4699 149773
rect 4389 140959 4699 149745
rect 4389 140931 4437 140959
rect 4465 140931 4499 140959
rect 4527 140931 4561 140959
rect 4589 140931 4623 140959
rect 4651 140931 4699 140959
rect 4389 140897 4699 140931
rect 4389 140869 4437 140897
rect 4465 140869 4499 140897
rect 4527 140869 4561 140897
rect 4589 140869 4623 140897
rect 4651 140869 4699 140897
rect 4389 140835 4699 140869
rect 4389 140807 4437 140835
rect 4465 140807 4499 140835
rect 4527 140807 4561 140835
rect 4589 140807 4623 140835
rect 4651 140807 4699 140835
rect 4389 140773 4699 140807
rect 4389 140745 4437 140773
rect 4465 140745 4499 140773
rect 4527 140745 4561 140773
rect 4589 140745 4623 140773
rect 4651 140745 4699 140773
rect 4389 131959 4699 140745
rect 4389 131931 4437 131959
rect 4465 131931 4499 131959
rect 4527 131931 4561 131959
rect 4589 131931 4623 131959
rect 4651 131931 4699 131959
rect 4389 131897 4699 131931
rect 4389 131869 4437 131897
rect 4465 131869 4499 131897
rect 4527 131869 4561 131897
rect 4589 131869 4623 131897
rect 4651 131869 4699 131897
rect 4389 131835 4699 131869
rect 4389 131807 4437 131835
rect 4465 131807 4499 131835
rect 4527 131807 4561 131835
rect 4589 131807 4623 131835
rect 4651 131807 4699 131835
rect 4389 131773 4699 131807
rect 4389 131745 4437 131773
rect 4465 131745 4499 131773
rect 4527 131745 4561 131773
rect 4589 131745 4623 131773
rect 4651 131745 4699 131773
rect 4389 122959 4699 131745
rect 4389 122931 4437 122959
rect 4465 122931 4499 122959
rect 4527 122931 4561 122959
rect 4589 122931 4623 122959
rect 4651 122931 4699 122959
rect 4389 122897 4699 122931
rect 4389 122869 4437 122897
rect 4465 122869 4499 122897
rect 4527 122869 4561 122897
rect 4589 122869 4623 122897
rect 4651 122869 4699 122897
rect 4389 122835 4699 122869
rect 4389 122807 4437 122835
rect 4465 122807 4499 122835
rect 4527 122807 4561 122835
rect 4589 122807 4623 122835
rect 4651 122807 4699 122835
rect 4389 122773 4699 122807
rect 4389 122745 4437 122773
rect 4465 122745 4499 122773
rect 4527 122745 4561 122773
rect 4589 122745 4623 122773
rect 4651 122745 4699 122773
rect 4389 113959 4699 122745
rect 4389 113931 4437 113959
rect 4465 113931 4499 113959
rect 4527 113931 4561 113959
rect 4589 113931 4623 113959
rect 4651 113931 4699 113959
rect 4389 113897 4699 113931
rect 4389 113869 4437 113897
rect 4465 113869 4499 113897
rect 4527 113869 4561 113897
rect 4589 113869 4623 113897
rect 4651 113869 4699 113897
rect 4389 113835 4699 113869
rect 4389 113807 4437 113835
rect 4465 113807 4499 113835
rect 4527 113807 4561 113835
rect 4589 113807 4623 113835
rect 4651 113807 4699 113835
rect 4389 113773 4699 113807
rect 4389 113745 4437 113773
rect 4465 113745 4499 113773
rect 4527 113745 4561 113773
rect 4589 113745 4623 113773
rect 4651 113745 4699 113773
rect 4389 104959 4699 113745
rect 4389 104931 4437 104959
rect 4465 104931 4499 104959
rect 4527 104931 4561 104959
rect 4589 104931 4623 104959
rect 4651 104931 4699 104959
rect 4389 104897 4699 104931
rect 4389 104869 4437 104897
rect 4465 104869 4499 104897
rect 4527 104869 4561 104897
rect 4589 104869 4623 104897
rect 4651 104869 4699 104897
rect 4389 104835 4699 104869
rect 4389 104807 4437 104835
rect 4465 104807 4499 104835
rect 4527 104807 4561 104835
rect 4589 104807 4623 104835
rect 4651 104807 4699 104835
rect 4389 104773 4699 104807
rect 4389 104745 4437 104773
rect 4465 104745 4499 104773
rect 4527 104745 4561 104773
rect 4589 104745 4623 104773
rect 4651 104745 4699 104773
rect 4389 95959 4699 104745
rect 4389 95931 4437 95959
rect 4465 95931 4499 95959
rect 4527 95931 4561 95959
rect 4589 95931 4623 95959
rect 4651 95931 4699 95959
rect 4389 95897 4699 95931
rect 4389 95869 4437 95897
rect 4465 95869 4499 95897
rect 4527 95869 4561 95897
rect 4589 95869 4623 95897
rect 4651 95869 4699 95897
rect 4389 95835 4699 95869
rect 4389 95807 4437 95835
rect 4465 95807 4499 95835
rect 4527 95807 4561 95835
rect 4589 95807 4623 95835
rect 4651 95807 4699 95835
rect 4389 95773 4699 95807
rect 4389 95745 4437 95773
rect 4465 95745 4499 95773
rect 4527 95745 4561 95773
rect 4589 95745 4623 95773
rect 4651 95745 4699 95773
rect 4389 86959 4699 95745
rect 4389 86931 4437 86959
rect 4465 86931 4499 86959
rect 4527 86931 4561 86959
rect 4589 86931 4623 86959
rect 4651 86931 4699 86959
rect 4389 86897 4699 86931
rect 4389 86869 4437 86897
rect 4465 86869 4499 86897
rect 4527 86869 4561 86897
rect 4589 86869 4623 86897
rect 4651 86869 4699 86897
rect 4389 86835 4699 86869
rect 4389 86807 4437 86835
rect 4465 86807 4499 86835
rect 4527 86807 4561 86835
rect 4589 86807 4623 86835
rect 4651 86807 4699 86835
rect 4389 86773 4699 86807
rect 4389 86745 4437 86773
rect 4465 86745 4499 86773
rect 4527 86745 4561 86773
rect 4589 86745 4623 86773
rect 4651 86745 4699 86773
rect 4389 77959 4699 86745
rect 4389 77931 4437 77959
rect 4465 77931 4499 77959
rect 4527 77931 4561 77959
rect 4589 77931 4623 77959
rect 4651 77931 4699 77959
rect 4389 77897 4699 77931
rect 4389 77869 4437 77897
rect 4465 77869 4499 77897
rect 4527 77869 4561 77897
rect 4589 77869 4623 77897
rect 4651 77869 4699 77897
rect 4389 77835 4699 77869
rect 4389 77807 4437 77835
rect 4465 77807 4499 77835
rect 4527 77807 4561 77835
rect 4589 77807 4623 77835
rect 4651 77807 4699 77835
rect 4389 77773 4699 77807
rect 4389 77745 4437 77773
rect 4465 77745 4499 77773
rect 4527 77745 4561 77773
rect 4589 77745 4623 77773
rect 4651 77745 4699 77773
rect 4389 68959 4699 77745
rect 4389 68931 4437 68959
rect 4465 68931 4499 68959
rect 4527 68931 4561 68959
rect 4589 68931 4623 68959
rect 4651 68931 4699 68959
rect 4389 68897 4699 68931
rect 4389 68869 4437 68897
rect 4465 68869 4499 68897
rect 4527 68869 4561 68897
rect 4589 68869 4623 68897
rect 4651 68869 4699 68897
rect 4389 68835 4699 68869
rect 4389 68807 4437 68835
rect 4465 68807 4499 68835
rect 4527 68807 4561 68835
rect 4589 68807 4623 68835
rect 4651 68807 4699 68835
rect 4389 68773 4699 68807
rect 4389 68745 4437 68773
rect 4465 68745 4499 68773
rect 4527 68745 4561 68773
rect 4589 68745 4623 68773
rect 4651 68745 4699 68773
rect 4389 59959 4699 68745
rect 4389 59931 4437 59959
rect 4465 59931 4499 59959
rect 4527 59931 4561 59959
rect 4589 59931 4623 59959
rect 4651 59931 4699 59959
rect 4389 59897 4699 59931
rect 4389 59869 4437 59897
rect 4465 59869 4499 59897
rect 4527 59869 4561 59897
rect 4589 59869 4623 59897
rect 4651 59869 4699 59897
rect 4389 59835 4699 59869
rect 4389 59807 4437 59835
rect 4465 59807 4499 59835
rect 4527 59807 4561 59835
rect 4589 59807 4623 59835
rect 4651 59807 4699 59835
rect 4389 59773 4699 59807
rect 4389 59745 4437 59773
rect 4465 59745 4499 59773
rect 4527 59745 4561 59773
rect 4589 59745 4623 59773
rect 4651 59745 4699 59773
rect 4389 50959 4699 59745
rect 4389 50931 4437 50959
rect 4465 50931 4499 50959
rect 4527 50931 4561 50959
rect 4589 50931 4623 50959
rect 4651 50931 4699 50959
rect 4389 50897 4699 50931
rect 4389 50869 4437 50897
rect 4465 50869 4499 50897
rect 4527 50869 4561 50897
rect 4589 50869 4623 50897
rect 4651 50869 4699 50897
rect 4389 50835 4699 50869
rect 4389 50807 4437 50835
rect 4465 50807 4499 50835
rect 4527 50807 4561 50835
rect 4589 50807 4623 50835
rect 4651 50807 4699 50835
rect 4389 50773 4699 50807
rect 4389 50745 4437 50773
rect 4465 50745 4499 50773
rect 4527 50745 4561 50773
rect 4589 50745 4623 50773
rect 4651 50745 4699 50773
rect 4389 41959 4699 50745
rect 4389 41931 4437 41959
rect 4465 41931 4499 41959
rect 4527 41931 4561 41959
rect 4589 41931 4623 41959
rect 4651 41931 4699 41959
rect 4389 41897 4699 41931
rect 4389 41869 4437 41897
rect 4465 41869 4499 41897
rect 4527 41869 4561 41897
rect 4589 41869 4623 41897
rect 4651 41869 4699 41897
rect 4389 41835 4699 41869
rect 4389 41807 4437 41835
rect 4465 41807 4499 41835
rect 4527 41807 4561 41835
rect 4589 41807 4623 41835
rect 4651 41807 4699 41835
rect 4389 41773 4699 41807
rect 4389 41745 4437 41773
rect 4465 41745 4499 41773
rect 4527 41745 4561 41773
rect 4589 41745 4623 41773
rect 4651 41745 4699 41773
rect 4389 32959 4699 41745
rect 4389 32931 4437 32959
rect 4465 32931 4499 32959
rect 4527 32931 4561 32959
rect 4589 32931 4623 32959
rect 4651 32931 4699 32959
rect 4389 32897 4699 32931
rect 4389 32869 4437 32897
rect 4465 32869 4499 32897
rect 4527 32869 4561 32897
rect 4589 32869 4623 32897
rect 4651 32869 4699 32897
rect 4389 32835 4699 32869
rect 4389 32807 4437 32835
rect 4465 32807 4499 32835
rect 4527 32807 4561 32835
rect 4589 32807 4623 32835
rect 4651 32807 4699 32835
rect 4389 32773 4699 32807
rect 4389 32745 4437 32773
rect 4465 32745 4499 32773
rect 4527 32745 4561 32773
rect 4589 32745 4623 32773
rect 4651 32745 4699 32773
rect 4389 23959 4699 32745
rect 4389 23931 4437 23959
rect 4465 23931 4499 23959
rect 4527 23931 4561 23959
rect 4589 23931 4623 23959
rect 4651 23931 4699 23959
rect 4389 23897 4699 23931
rect 4389 23869 4437 23897
rect 4465 23869 4499 23897
rect 4527 23869 4561 23897
rect 4589 23869 4623 23897
rect 4651 23869 4699 23897
rect 4389 23835 4699 23869
rect 4389 23807 4437 23835
rect 4465 23807 4499 23835
rect 4527 23807 4561 23835
rect 4589 23807 4623 23835
rect 4651 23807 4699 23835
rect 4389 23773 4699 23807
rect 4389 23745 4437 23773
rect 4465 23745 4499 23773
rect 4527 23745 4561 23773
rect 4589 23745 4623 23773
rect 4651 23745 4699 23773
rect 4389 14959 4699 23745
rect 4389 14931 4437 14959
rect 4465 14931 4499 14959
rect 4527 14931 4561 14959
rect 4589 14931 4623 14959
rect 4651 14931 4699 14959
rect 4389 14897 4699 14931
rect 4389 14869 4437 14897
rect 4465 14869 4499 14897
rect 4527 14869 4561 14897
rect 4589 14869 4623 14897
rect 4651 14869 4699 14897
rect 4389 14835 4699 14869
rect 4389 14807 4437 14835
rect 4465 14807 4499 14835
rect 4527 14807 4561 14835
rect 4589 14807 4623 14835
rect 4651 14807 4699 14835
rect 4389 14773 4699 14807
rect 4389 14745 4437 14773
rect 4465 14745 4499 14773
rect 4527 14745 4561 14773
rect 4589 14745 4623 14773
rect 4651 14745 4699 14773
rect 4389 5959 4699 14745
rect 4389 5931 4437 5959
rect 4465 5931 4499 5959
rect 4527 5931 4561 5959
rect 4589 5931 4623 5959
rect 4651 5931 4699 5959
rect 4389 5897 4699 5931
rect 4389 5869 4437 5897
rect 4465 5869 4499 5897
rect 4527 5869 4561 5897
rect 4589 5869 4623 5897
rect 4651 5869 4699 5897
rect 4389 5835 4699 5869
rect 4389 5807 4437 5835
rect 4465 5807 4499 5835
rect 4527 5807 4561 5835
rect 4589 5807 4623 5835
rect 4651 5807 4699 5835
rect 4389 5773 4699 5807
rect 4389 5745 4437 5773
rect 4465 5745 4499 5773
rect 4527 5745 4561 5773
rect 4589 5745 4623 5773
rect 4651 5745 4699 5773
rect 4389 424 4699 5745
rect 4389 396 4437 424
rect 4465 396 4499 424
rect 4527 396 4561 424
rect 4589 396 4623 424
rect 4651 396 4699 424
rect 4389 362 4699 396
rect 4389 334 4437 362
rect 4465 334 4499 362
rect 4527 334 4561 362
rect 4589 334 4623 362
rect 4651 334 4699 362
rect 4389 300 4699 334
rect 4389 272 4437 300
rect 4465 272 4499 300
rect 4527 272 4561 300
rect 4589 272 4623 300
rect 4651 272 4699 300
rect 4389 238 4699 272
rect 4389 210 4437 238
rect 4465 210 4499 238
rect 4527 210 4561 238
rect 4589 210 4623 238
rect 4651 210 4699 238
rect 4389 162 4699 210
rect 11529 299190 11839 299718
rect 11529 299162 11577 299190
rect 11605 299162 11639 299190
rect 11667 299162 11701 299190
rect 11729 299162 11763 299190
rect 11791 299162 11839 299190
rect 11529 299128 11839 299162
rect 11529 299100 11577 299128
rect 11605 299100 11639 299128
rect 11667 299100 11701 299128
rect 11729 299100 11763 299128
rect 11791 299100 11839 299128
rect 11529 299066 11839 299100
rect 11529 299038 11577 299066
rect 11605 299038 11639 299066
rect 11667 299038 11701 299066
rect 11729 299038 11763 299066
rect 11791 299038 11839 299066
rect 11529 299004 11839 299038
rect 11529 298976 11577 299004
rect 11605 298976 11639 299004
rect 11667 298976 11701 299004
rect 11729 298976 11763 299004
rect 11791 298976 11839 299004
rect 11529 290959 11839 298976
rect 11529 290931 11577 290959
rect 11605 290931 11639 290959
rect 11667 290931 11701 290959
rect 11729 290931 11763 290959
rect 11791 290931 11839 290959
rect 11529 290897 11839 290931
rect 11529 290869 11577 290897
rect 11605 290869 11639 290897
rect 11667 290869 11701 290897
rect 11729 290869 11763 290897
rect 11791 290869 11839 290897
rect 11529 290835 11839 290869
rect 11529 290807 11577 290835
rect 11605 290807 11639 290835
rect 11667 290807 11701 290835
rect 11729 290807 11763 290835
rect 11791 290807 11839 290835
rect 11529 290773 11839 290807
rect 11529 290745 11577 290773
rect 11605 290745 11639 290773
rect 11667 290745 11701 290773
rect 11729 290745 11763 290773
rect 11791 290745 11839 290773
rect 11529 281959 11839 290745
rect 11529 281931 11577 281959
rect 11605 281931 11639 281959
rect 11667 281931 11701 281959
rect 11729 281931 11763 281959
rect 11791 281931 11839 281959
rect 11529 281897 11839 281931
rect 11529 281869 11577 281897
rect 11605 281869 11639 281897
rect 11667 281869 11701 281897
rect 11729 281869 11763 281897
rect 11791 281869 11839 281897
rect 11529 281835 11839 281869
rect 11529 281807 11577 281835
rect 11605 281807 11639 281835
rect 11667 281807 11701 281835
rect 11729 281807 11763 281835
rect 11791 281807 11839 281835
rect 11529 281773 11839 281807
rect 11529 281745 11577 281773
rect 11605 281745 11639 281773
rect 11667 281745 11701 281773
rect 11729 281745 11763 281773
rect 11791 281745 11839 281773
rect 11529 272959 11839 281745
rect 11529 272931 11577 272959
rect 11605 272931 11639 272959
rect 11667 272931 11701 272959
rect 11729 272931 11763 272959
rect 11791 272931 11839 272959
rect 11529 272897 11839 272931
rect 11529 272869 11577 272897
rect 11605 272869 11639 272897
rect 11667 272869 11701 272897
rect 11729 272869 11763 272897
rect 11791 272869 11839 272897
rect 11529 272835 11839 272869
rect 11529 272807 11577 272835
rect 11605 272807 11639 272835
rect 11667 272807 11701 272835
rect 11729 272807 11763 272835
rect 11791 272807 11839 272835
rect 11529 272773 11839 272807
rect 11529 272745 11577 272773
rect 11605 272745 11639 272773
rect 11667 272745 11701 272773
rect 11729 272745 11763 272773
rect 11791 272745 11839 272773
rect 11529 263959 11839 272745
rect 11529 263931 11577 263959
rect 11605 263931 11639 263959
rect 11667 263931 11701 263959
rect 11729 263931 11763 263959
rect 11791 263931 11839 263959
rect 11529 263897 11839 263931
rect 11529 263869 11577 263897
rect 11605 263869 11639 263897
rect 11667 263869 11701 263897
rect 11729 263869 11763 263897
rect 11791 263869 11839 263897
rect 11529 263835 11839 263869
rect 11529 263807 11577 263835
rect 11605 263807 11639 263835
rect 11667 263807 11701 263835
rect 11729 263807 11763 263835
rect 11791 263807 11839 263835
rect 11529 263773 11839 263807
rect 11529 263745 11577 263773
rect 11605 263745 11639 263773
rect 11667 263745 11701 263773
rect 11729 263745 11763 263773
rect 11791 263745 11839 263773
rect 11529 254959 11839 263745
rect 11529 254931 11577 254959
rect 11605 254931 11639 254959
rect 11667 254931 11701 254959
rect 11729 254931 11763 254959
rect 11791 254931 11839 254959
rect 11529 254897 11839 254931
rect 11529 254869 11577 254897
rect 11605 254869 11639 254897
rect 11667 254869 11701 254897
rect 11729 254869 11763 254897
rect 11791 254869 11839 254897
rect 11529 254835 11839 254869
rect 11529 254807 11577 254835
rect 11605 254807 11639 254835
rect 11667 254807 11701 254835
rect 11729 254807 11763 254835
rect 11791 254807 11839 254835
rect 11529 254773 11839 254807
rect 11529 254745 11577 254773
rect 11605 254745 11639 254773
rect 11667 254745 11701 254773
rect 11729 254745 11763 254773
rect 11791 254745 11839 254773
rect 11529 245959 11839 254745
rect 11529 245931 11577 245959
rect 11605 245931 11639 245959
rect 11667 245931 11701 245959
rect 11729 245931 11763 245959
rect 11791 245931 11839 245959
rect 11529 245897 11839 245931
rect 11529 245869 11577 245897
rect 11605 245869 11639 245897
rect 11667 245869 11701 245897
rect 11729 245869 11763 245897
rect 11791 245869 11839 245897
rect 11529 245835 11839 245869
rect 11529 245807 11577 245835
rect 11605 245807 11639 245835
rect 11667 245807 11701 245835
rect 11729 245807 11763 245835
rect 11791 245807 11839 245835
rect 11529 245773 11839 245807
rect 11529 245745 11577 245773
rect 11605 245745 11639 245773
rect 11667 245745 11701 245773
rect 11729 245745 11763 245773
rect 11791 245745 11839 245773
rect 11529 236959 11839 245745
rect 11529 236931 11577 236959
rect 11605 236931 11639 236959
rect 11667 236931 11701 236959
rect 11729 236931 11763 236959
rect 11791 236931 11839 236959
rect 11529 236897 11839 236931
rect 11529 236869 11577 236897
rect 11605 236869 11639 236897
rect 11667 236869 11701 236897
rect 11729 236869 11763 236897
rect 11791 236869 11839 236897
rect 11529 236835 11839 236869
rect 11529 236807 11577 236835
rect 11605 236807 11639 236835
rect 11667 236807 11701 236835
rect 11729 236807 11763 236835
rect 11791 236807 11839 236835
rect 11529 236773 11839 236807
rect 11529 236745 11577 236773
rect 11605 236745 11639 236773
rect 11667 236745 11701 236773
rect 11729 236745 11763 236773
rect 11791 236745 11839 236773
rect 11529 227959 11839 236745
rect 11529 227931 11577 227959
rect 11605 227931 11639 227959
rect 11667 227931 11701 227959
rect 11729 227931 11763 227959
rect 11791 227931 11839 227959
rect 11529 227897 11839 227931
rect 11529 227869 11577 227897
rect 11605 227869 11639 227897
rect 11667 227869 11701 227897
rect 11729 227869 11763 227897
rect 11791 227869 11839 227897
rect 11529 227835 11839 227869
rect 11529 227807 11577 227835
rect 11605 227807 11639 227835
rect 11667 227807 11701 227835
rect 11729 227807 11763 227835
rect 11791 227807 11839 227835
rect 11529 227773 11839 227807
rect 11529 227745 11577 227773
rect 11605 227745 11639 227773
rect 11667 227745 11701 227773
rect 11729 227745 11763 227773
rect 11791 227745 11839 227773
rect 11529 218959 11839 227745
rect 11529 218931 11577 218959
rect 11605 218931 11639 218959
rect 11667 218931 11701 218959
rect 11729 218931 11763 218959
rect 11791 218931 11839 218959
rect 11529 218897 11839 218931
rect 11529 218869 11577 218897
rect 11605 218869 11639 218897
rect 11667 218869 11701 218897
rect 11729 218869 11763 218897
rect 11791 218869 11839 218897
rect 11529 218835 11839 218869
rect 11529 218807 11577 218835
rect 11605 218807 11639 218835
rect 11667 218807 11701 218835
rect 11729 218807 11763 218835
rect 11791 218807 11839 218835
rect 11529 218773 11839 218807
rect 11529 218745 11577 218773
rect 11605 218745 11639 218773
rect 11667 218745 11701 218773
rect 11729 218745 11763 218773
rect 11791 218745 11839 218773
rect 11529 209959 11839 218745
rect 11529 209931 11577 209959
rect 11605 209931 11639 209959
rect 11667 209931 11701 209959
rect 11729 209931 11763 209959
rect 11791 209931 11839 209959
rect 11529 209897 11839 209931
rect 11529 209869 11577 209897
rect 11605 209869 11639 209897
rect 11667 209869 11701 209897
rect 11729 209869 11763 209897
rect 11791 209869 11839 209897
rect 11529 209835 11839 209869
rect 11529 209807 11577 209835
rect 11605 209807 11639 209835
rect 11667 209807 11701 209835
rect 11729 209807 11763 209835
rect 11791 209807 11839 209835
rect 11529 209773 11839 209807
rect 11529 209745 11577 209773
rect 11605 209745 11639 209773
rect 11667 209745 11701 209773
rect 11729 209745 11763 209773
rect 11791 209745 11839 209773
rect 11529 200959 11839 209745
rect 11529 200931 11577 200959
rect 11605 200931 11639 200959
rect 11667 200931 11701 200959
rect 11729 200931 11763 200959
rect 11791 200931 11839 200959
rect 11529 200897 11839 200931
rect 11529 200869 11577 200897
rect 11605 200869 11639 200897
rect 11667 200869 11701 200897
rect 11729 200869 11763 200897
rect 11791 200869 11839 200897
rect 11529 200835 11839 200869
rect 11529 200807 11577 200835
rect 11605 200807 11639 200835
rect 11667 200807 11701 200835
rect 11729 200807 11763 200835
rect 11791 200807 11839 200835
rect 11529 200773 11839 200807
rect 11529 200745 11577 200773
rect 11605 200745 11639 200773
rect 11667 200745 11701 200773
rect 11729 200745 11763 200773
rect 11791 200745 11839 200773
rect 11529 191959 11839 200745
rect 11529 191931 11577 191959
rect 11605 191931 11639 191959
rect 11667 191931 11701 191959
rect 11729 191931 11763 191959
rect 11791 191931 11839 191959
rect 11529 191897 11839 191931
rect 11529 191869 11577 191897
rect 11605 191869 11639 191897
rect 11667 191869 11701 191897
rect 11729 191869 11763 191897
rect 11791 191869 11839 191897
rect 11529 191835 11839 191869
rect 11529 191807 11577 191835
rect 11605 191807 11639 191835
rect 11667 191807 11701 191835
rect 11729 191807 11763 191835
rect 11791 191807 11839 191835
rect 11529 191773 11839 191807
rect 11529 191745 11577 191773
rect 11605 191745 11639 191773
rect 11667 191745 11701 191773
rect 11729 191745 11763 191773
rect 11791 191745 11839 191773
rect 11529 182959 11839 191745
rect 11529 182931 11577 182959
rect 11605 182931 11639 182959
rect 11667 182931 11701 182959
rect 11729 182931 11763 182959
rect 11791 182931 11839 182959
rect 11529 182897 11839 182931
rect 11529 182869 11577 182897
rect 11605 182869 11639 182897
rect 11667 182869 11701 182897
rect 11729 182869 11763 182897
rect 11791 182869 11839 182897
rect 11529 182835 11839 182869
rect 11529 182807 11577 182835
rect 11605 182807 11639 182835
rect 11667 182807 11701 182835
rect 11729 182807 11763 182835
rect 11791 182807 11839 182835
rect 11529 182773 11839 182807
rect 11529 182745 11577 182773
rect 11605 182745 11639 182773
rect 11667 182745 11701 182773
rect 11729 182745 11763 182773
rect 11791 182745 11839 182773
rect 11529 173959 11839 182745
rect 11529 173931 11577 173959
rect 11605 173931 11639 173959
rect 11667 173931 11701 173959
rect 11729 173931 11763 173959
rect 11791 173931 11839 173959
rect 11529 173897 11839 173931
rect 11529 173869 11577 173897
rect 11605 173869 11639 173897
rect 11667 173869 11701 173897
rect 11729 173869 11763 173897
rect 11791 173869 11839 173897
rect 11529 173835 11839 173869
rect 11529 173807 11577 173835
rect 11605 173807 11639 173835
rect 11667 173807 11701 173835
rect 11729 173807 11763 173835
rect 11791 173807 11839 173835
rect 11529 173773 11839 173807
rect 11529 173745 11577 173773
rect 11605 173745 11639 173773
rect 11667 173745 11701 173773
rect 11729 173745 11763 173773
rect 11791 173745 11839 173773
rect 11529 164959 11839 173745
rect 11529 164931 11577 164959
rect 11605 164931 11639 164959
rect 11667 164931 11701 164959
rect 11729 164931 11763 164959
rect 11791 164931 11839 164959
rect 11529 164897 11839 164931
rect 11529 164869 11577 164897
rect 11605 164869 11639 164897
rect 11667 164869 11701 164897
rect 11729 164869 11763 164897
rect 11791 164869 11839 164897
rect 11529 164835 11839 164869
rect 11529 164807 11577 164835
rect 11605 164807 11639 164835
rect 11667 164807 11701 164835
rect 11729 164807 11763 164835
rect 11791 164807 11839 164835
rect 11529 164773 11839 164807
rect 11529 164745 11577 164773
rect 11605 164745 11639 164773
rect 11667 164745 11701 164773
rect 11729 164745 11763 164773
rect 11791 164745 11839 164773
rect 11529 155959 11839 164745
rect 11529 155931 11577 155959
rect 11605 155931 11639 155959
rect 11667 155931 11701 155959
rect 11729 155931 11763 155959
rect 11791 155931 11839 155959
rect 11529 155897 11839 155931
rect 11529 155869 11577 155897
rect 11605 155869 11639 155897
rect 11667 155869 11701 155897
rect 11729 155869 11763 155897
rect 11791 155869 11839 155897
rect 11529 155835 11839 155869
rect 11529 155807 11577 155835
rect 11605 155807 11639 155835
rect 11667 155807 11701 155835
rect 11729 155807 11763 155835
rect 11791 155807 11839 155835
rect 11529 155773 11839 155807
rect 11529 155745 11577 155773
rect 11605 155745 11639 155773
rect 11667 155745 11701 155773
rect 11729 155745 11763 155773
rect 11791 155745 11839 155773
rect 11529 146959 11839 155745
rect 11529 146931 11577 146959
rect 11605 146931 11639 146959
rect 11667 146931 11701 146959
rect 11729 146931 11763 146959
rect 11791 146931 11839 146959
rect 11529 146897 11839 146931
rect 11529 146869 11577 146897
rect 11605 146869 11639 146897
rect 11667 146869 11701 146897
rect 11729 146869 11763 146897
rect 11791 146869 11839 146897
rect 11529 146835 11839 146869
rect 11529 146807 11577 146835
rect 11605 146807 11639 146835
rect 11667 146807 11701 146835
rect 11729 146807 11763 146835
rect 11791 146807 11839 146835
rect 11529 146773 11839 146807
rect 11529 146745 11577 146773
rect 11605 146745 11639 146773
rect 11667 146745 11701 146773
rect 11729 146745 11763 146773
rect 11791 146745 11839 146773
rect 11529 137959 11839 146745
rect 11529 137931 11577 137959
rect 11605 137931 11639 137959
rect 11667 137931 11701 137959
rect 11729 137931 11763 137959
rect 11791 137931 11839 137959
rect 11529 137897 11839 137931
rect 11529 137869 11577 137897
rect 11605 137869 11639 137897
rect 11667 137869 11701 137897
rect 11729 137869 11763 137897
rect 11791 137869 11839 137897
rect 11529 137835 11839 137869
rect 11529 137807 11577 137835
rect 11605 137807 11639 137835
rect 11667 137807 11701 137835
rect 11729 137807 11763 137835
rect 11791 137807 11839 137835
rect 11529 137773 11839 137807
rect 11529 137745 11577 137773
rect 11605 137745 11639 137773
rect 11667 137745 11701 137773
rect 11729 137745 11763 137773
rect 11791 137745 11839 137773
rect 11529 128959 11839 137745
rect 11529 128931 11577 128959
rect 11605 128931 11639 128959
rect 11667 128931 11701 128959
rect 11729 128931 11763 128959
rect 11791 128931 11839 128959
rect 11529 128897 11839 128931
rect 11529 128869 11577 128897
rect 11605 128869 11639 128897
rect 11667 128869 11701 128897
rect 11729 128869 11763 128897
rect 11791 128869 11839 128897
rect 11529 128835 11839 128869
rect 11529 128807 11577 128835
rect 11605 128807 11639 128835
rect 11667 128807 11701 128835
rect 11729 128807 11763 128835
rect 11791 128807 11839 128835
rect 11529 128773 11839 128807
rect 11529 128745 11577 128773
rect 11605 128745 11639 128773
rect 11667 128745 11701 128773
rect 11729 128745 11763 128773
rect 11791 128745 11839 128773
rect 11529 119959 11839 128745
rect 11529 119931 11577 119959
rect 11605 119931 11639 119959
rect 11667 119931 11701 119959
rect 11729 119931 11763 119959
rect 11791 119931 11839 119959
rect 11529 119897 11839 119931
rect 11529 119869 11577 119897
rect 11605 119869 11639 119897
rect 11667 119869 11701 119897
rect 11729 119869 11763 119897
rect 11791 119869 11839 119897
rect 11529 119835 11839 119869
rect 11529 119807 11577 119835
rect 11605 119807 11639 119835
rect 11667 119807 11701 119835
rect 11729 119807 11763 119835
rect 11791 119807 11839 119835
rect 11529 119773 11839 119807
rect 11529 119745 11577 119773
rect 11605 119745 11639 119773
rect 11667 119745 11701 119773
rect 11729 119745 11763 119773
rect 11791 119745 11839 119773
rect 11529 110959 11839 119745
rect 11529 110931 11577 110959
rect 11605 110931 11639 110959
rect 11667 110931 11701 110959
rect 11729 110931 11763 110959
rect 11791 110931 11839 110959
rect 11529 110897 11839 110931
rect 11529 110869 11577 110897
rect 11605 110869 11639 110897
rect 11667 110869 11701 110897
rect 11729 110869 11763 110897
rect 11791 110869 11839 110897
rect 11529 110835 11839 110869
rect 11529 110807 11577 110835
rect 11605 110807 11639 110835
rect 11667 110807 11701 110835
rect 11729 110807 11763 110835
rect 11791 110807 11839 110835
rect 11529 110773 11839 110807
rect 11529 110745 11577 110773
rect 11605 110745 11639 110773
rect 11667 110745 11701 110773
rect 11729 110745 11763 110773
rect 11791 110745 11839 110773
rect 11529 101959 11839 110745
rect 11529 101931 11577 101959
rect 11605 101931 11639 101959
rect 11667 101931 11701 101959
rect 11729 101931 11763 101959
rect 11791 101931 11839 101959
rect 11529 101897 11839 101931
rect 11529 101869 11577 101897
rect 11605 101869 11639 101897
rect 11667 101869 11701 101897
rect 11729 101869 11763 101897
rect 11791 101869 11839 101897
rect 11529 101835 11839 101869
rect 11529 101807 11577 101835
rect 11605 101807 11639 101835
rect 11667 101807 11701 101835
rect 11729 101807 11763 101835
rect 11791 101807 11839 101835
rect 11529 101773 11839 101807
rect 11529 101745 11577 101773
rect 11605 101745 11639 101773
rect 11667 101745 11701 101773
rect 11729 101745 11763 101773
rect 11791 101745 11839 101773
rect 11529 92959 11839 101745
rect 11529 92931 11577 92959
rect 11605 92931 11639 92959
rect 11667 92931 11701 92959
rect 11729 92931 11763 92959
rect 11791 92931 11839 92959
rect 11529 92897 11839 92931
rect 11529 92869 11577 92897
rect 11605 92869 11639 92897
rect 11667 92869 11701 92897
rect 11729 92869 11763 92897
rect 11791 92869 11839 92897
rect 11529 92835 11839 92869
rect 11529 92807 11577 92835
rect 11605 92807 11639 92835
rect 11667 92807 11701 92835
rect 11729 92807 11763 92835
rect 11791 92807 11839 92835
rect 11529 92773 11839 92807
rect 11529 92745 11577 92773
rect 11605 92745 11639 92773
rect 11667 92745 11701 92773
rect 11729 92745 11763 92773
rect 11791 92745 11839 92773
rect 11529 83959 11839 92745
rect 11529 83931 11577 83959
rect 11605 83931 11639 83959
rect 11667 83931 11701 83959
rect 11729 83931 11763 83959
rect 11791 83931 11839 83959
rect 11529 83897 11839 83931
rect 11529 83869 11577 83897
rect 11605 83869 11639 83897
rect 11667 83869 11701 83897
rect 11729 83869 11763 83897
rect 11791 83869 11839 83897
rect 11529 83835 11839 83869
rect 11529 83807 11577 83835
rect 11605 83807 11639 83835
rect 11667 83807 11701 83835
rect 11729 83807 11763 83835
rect 11791 83807 11839 83835
rect 11529 83773 11839 83807
rect 11529 83745 11577 83773
rect 11605 83745 11639 83773
rect 11667 83745 11701 83773
rect 11729 83745 11763 83773
rect 11791 83745 11839 83773
rect 11529 74959 11839 83745
rect 11529 74931 11577 74959
rect 11605 74931 11639 74959
rect 11667 74931 11701 74959
rect 11729 74931 11763 74959
rect 11791 74931 11839 74959
rect 11529 74897 11839 74931
rect 11529 74869 11577 74897
rect 11605 74869 11639 74897
rect 11667 74869 11701 74897
rect 11729 74869 11763 74897
rect 11791 74869 11839 74897
rect 11529 74835 11839 74869
rect 11529 74807 11577 74835
rect 11605 74807 11639 74835
rect 11667 74807 11701 74835
rect 11729 74807 11763 74835
rect 11791 74807 11839 74835
rect 11529 74773 11839 74807
rect 11529 74745 11577 74773
rect 11605 74745 11639 74773
rect 11667 74745 11701 74773
rect 11729 74745 11763 74773
rect 11791 74745 11839 74773
rect 11529 65959 11839 74745
rect 11529 65931 11577 65959
rect 11605 65931 11639 65959
rect 11667 65931 11701 65959
rect 11729 65931 11763 65959
rect 11791 65931 11839 65959
rect 11529 65897 11839 65931
rect 11529 65869 11577 65897
rect 11605 65869 11639 65897
rect 11667 65869 11701 65897
rect 11729 65869 11763 65897
rect 11791 65869 11839 65897
rect 11529 65835 11839 65869
rect 11529 65807 11577 65835
rect 11605 65807 11639 65835
rect 11667 65807 11701 65835
rect 11729 65807 11763 65835
rect 11791 65807 11839 65835
rect 11529 65773 11839 65807
rect 11529 65745 11577 65773
rect 11605 65745 11639 65773
rect 11667 65745 11701 65773
rect 11729 65745 11763 65773
rect 11791 65745 11839 65773
rect 11529 56959 11839 65745
rect 11529 56931 11577 56959
rect 11605 56931 11639 56959
rect 11667 56931 11701 56959
rect 11729 56931 11763 56959
rect 11791 56931 11839 56959
rect 11529 56897 11839 56931
rect 11529 56869 11577 56897
rect 11605 56869 11639 56897
rect 11667 56869 11701 56897
rect 11729 56869 11763 56897
rect 11791 56869 11839 56897
rect 11529 56835 11839 56869
rect 11529 56807 11577 56835
rect 11605 56807 11639 56835
rect 11667 56807 11701 56835
rect 11729 56807 11763 56835
rect 11791 56807 11839 56835
rect 11529 56773 11839 56807
rect 11529 56745 11577 56773
rect 11605 56745 11639 56773
rect 11667 56745 11701 56773
rect 11729 56745 11763 56773
rect 11791 56745 11839 56773
rect 11529 47959 11839 56745
rect 11529 47931 11577 47959
rect 11605 47931 11639 47959
rect 11667 47931 11701 47959
rect 11729 47931 11763 47959
rect 11791 47931 11839 47959
rect 11529 47897 11839 47931
rect 11529 47869 11577 47897
rect 11605 47869 11639 47897
rect 11667 47869 11701 47897
rect 11729 47869 11763 47897
rect 11791 47869 11839 47897
rect 11529 47835 11839 47869
rect 11529 47807 11577 47835
rect 11605 47807 11639 47835
rect 11667 47807 11701 47835
rect 11729 47807 11763 47835
rect 11791 47807 11839 47835
rect 11529 47773 11839 47807
rect 11529 47745 11577 47773
rect 11605 47745 11639 47773
rect 11667 47745 11701 47773
rect 11729 47745 11763 47773
rect 11791 47745 11839 47773
rect 11529 38959 11839 47745
rect 11529 38931 11577 38959
rect 11605 38931 11639 38959
rect 11667 38931 11701 38959
rect 11729 38931 11763 38959
rect 11791 38931 11839 38959
rect 11529 38897 11839 38931
rect 11529 38869 11577 38897
rect 11605 38869 11639 38897
rect 11667 38869 11701 38897
rect 11729 38869 11763 38897
rect 11791 38869 11839 38897
rect 11529 38835 11839 38869
rect 11529 38807 11577 38835
rect 11605 38807 11639 38835
rect 11667 38807 11701 38835
rect 11729 38807 11763 38835
rect 11791 38807 11839 38835
rect 11529 38773 11839 38807
rect 11529 38745 11577 38773
rect 11605 38745 11639 38773
rect 11667 38745 11701 38773
rect 11729 38745 11763 38773
rect 11791 38745 11839 38773
rect 11529 29959 11839 38745
rect 11529 29931 11577 29959
rect 11605 29931 11639 29959
rect 11667 29931 11701 29959
rect 11729 29931 11763 29959
rect 11791 29931 11839 29959
rect 11529 29897 11839 29931
rect 11529 29869 11577 29897
rect 11605 29869 11639 29897
rect 11667 29869 11701 29897
rect 11729 29869 11763 29897
rect 11791 29869 11839 29897
rect 11529 29835 11839 29869
rect 11529 29807 11577 29835
rect 11605 29807 11639 29835
rect 11667 29807 11701 29835
rect 11729 29807 11763 29835
rect 11791 29807 11839 29835
rect 11529 29773 11839 29807
rect 11529 29745 11577 29773
rect 11605 29745 11639 29773
rect 11667 29745 11701 29773
rect 11729 29745 11763 29773
rect 11791 29745 11839 29773
rect 11529 20959 11839 29745
rect 11529 20931 11577 20959
rect 11605 20931 11639 20959
rect 11667 20931 11701 20959
rect 11729 20931 11763 20959
rect 11791 20931 11839 20959
rect 11529 20897 11839 20931
rect 11529 20869 11577 20897
rect 11605 20869 11639 20897
rect 11667 20869 11701 20897
rect 11729 20869 11763 20897
rect 11791 20869 11839 20897
rect 11529 20835 11839 20869
rect 11529 20807 11577 20835
rect 11605 20807 11639 20835
rect 11667 20807 11701 20835
rect 11729 20807 11763 20835
rect 11791 20807 11839 20835
rect 11529 20773 11839 20807
rect 11529 20745 11577 20773
rect 11605 20745 11639 20773
rect 11667 20745 11701 20773
rect 11729 20745 11763 20773
rect 11791 20745 11839 20773
rect 11529 11959 11839 20745
rect 11529 11931 11577 11959
rect 11605 11931 11639 11959
rect 11667 11931 11701 11959
rect 11729 11931 11763 11959
rect 11791 11931 11839 11959
rect 11529 11897 11839 11931
rect 11529 11869 11577 11897
rect 11605 11869 11639 11897
rect 11667 11869 11701 11897
rect 11729 11869 11763 11897
rect 11791 11869 11839 11897
rect 11529 11835 11839 11869
rect 11529 11807 11577 11835
rect 11605 11807 11639 11835
rect 11667 11807 11701 11835
rect 11729 11807 11763 11835
rect 11791 11807 11839 11835
rect 11529 11773 11839 11807
rect 11529 11745 11577 11773
rect 11605 11745 11639 11773
rect 11667 11745 11701 11773
rect 11729 11745 11763 11773
rect 11791 11745 11839 11773
rect 11529 2959 11839 11745
rect 11529 2931 11577 2959
rect 11605 2931 11639 2959
rect 11667 2931 11701 2959
rect 11729 2931 11763 2959
rect 11791 2931 11839 2959
rect 11529 2897 11839 2931
rect 11529 2869 11577 2897
rect 11605 2869 11639 2897
rect 11667 2869 11701 2897
rect 11729 2869 11763 2897
rect 11791 2869 11839 2897
rect 11529 2835 11839 2869
rect 11529 2807 11577 2835
rect 11605 2807 11639 2835
rect 11667 2807 11701 2835
rect 11729 2807 11763 2835
rect 11791 2807 11839 2835
rect 11529 2773 11839 2807
rect 11529 2745 11577 2773
rect 11605 2745 11639 2773
rect 11667 2745 11701 2773
rect 11729 2745 11763 2773
rect 11791 2745 11839 2773
rect 11529 904 11839 2745
rect 11529 876 11577 904
rect 11605 876 11639 904
rect 11667 876 11701 904
rect 11729 876 11763 904
rect 11791 876 11839 904
rect 11529 842 11839 876
rect 11529 814 11577 842
rect 11605 814 11639 842
rect 11667 814 11701 842
rect 11729 814 11763 842
rect 11791 814 11839 842
rect 11529 780 11839 814
rect 11529 752 11577 780
rect 11605 752 11639 780
rect 11667 752 11701 780
rect 11729 752 11763 780
rect 11791 752 11839 780
rect 11529 718 11839 752
rect 11529 690 11577 718
rect 11605 690 11639 718
rect 11667 690 11701 718
rect 11729 690 11763 718
rect 11791 690 11839 718
rect 11529 162 11839 690
rect 13389 299670 13699 299718
rect 13389 299642 13437 299670
rect 13465 299642 13499 299670
rect 13527 299642 13561 299670
rect 13589 299642 13623 299670
rect 13651 299642 13699 299670
rect 13389 299608 13699 299642
rect 13389 299580 13437 299608
rect 13465 299580 13499 299608
rect 13527 299580 13561 299608
rect 13589 299580 13623 299608
rect 13651 299580 13699 299608
rect 13389 299546 13699 299580
rect 13389 299518 13437 299546
rect 13465 299518 13499 299546
rect 13527 299518 13561 299546
rect 13589 299518 13623 299546
rect 13651 299518 13699 299546
rect 13389 299484 13699 299518
rect 13389 299456 13437 299484
rect 13465 299456 13499 299484
rect 13527 299456 13561 299484
rect 13589 299456 13623 299484
rect 13651 299456 13699 299484
rect 13389 293959 13699 299456
rect 13389 293931 13437 293959
rect 13465 293931 13499 293959
rect 13527 293931 13561 293959
rect 13589 293931 13623 293959
rect 13651 293931 13699 293959
rect 13389 293897 13699 293931
rect 13389 293869 13437 293897
rect 13465 293869 13499 293897
rect 13527 293869 13561 293897
rect 13589 293869 13623 293897
rect 13651 293869 13699 293897
rect 13389 293835 13699 293869
rect 13389 293807 13437 293835
rect 13465 293807 13499 293835
rect 13527 293807 13561 293835
rect 13589 293807 13623 293835
rect 13651 293807 13699 293835
rect 13389 293773 13699 293807
rect 13389 293745 13437 293773
rect 13465 293745 13499 293773
rect 13527 293745 13561 293773
rect 13589 293745 13623 293773
rect 13651 293745 13699 293773
rect 13389 284959 13699 293745
rect 13389 284931 13437 284959
rect 13465 284931 13499 284959
rect 13527 284931 13561 284959
rect 13589 284931 13623 284959
rect 13651 284931 13699 284959
rect 13389 284897 13699 284931
rect 13389 284869 13437 284897
rect 13465 284869 13499 284897
rect 13527 284869 13561 284897
rect 13589 284869 13623 284897
rect 13651 284869 13699 284897
rect 13389 284835 13699 284869
rect 13389 284807 13437 284835
rect 13465 284807 13499 284835
rect 13527 284807 13561 284835
rect 13589 284807 13623 284835
rect 13651 284807 13699 284835
rect 13389 284773 13699 284807
rect 13389 284745 13437 284773
rect 13465 284745 13499 284773
rect 13527 284745 13561 284773
rect 13589 284745 13623 284773
rect 13651 284745 13699 284773
rect 13389 275959 13699 284745
rect 13389 275931 13437 275959
rect 13465 275931 13499 275959
rect 13527 275931 13561 275959
rect 13589 275931 13623 275959
rect 13651 275931 13699 275959
rect 13389 275897 13699 275931
rect 13389 275869 13437 275897
rect 13465 275869 13499 275897
rect 13527 275869 13561 275897
rect 13589 275869 13623 275897
rect 13651 275869 13699 275897
rect 13389 275835 13699 275869
rect 13389 275807 13437 275835
rect 13465 275807 13499 275835
rect 13527 275807 13561 275835
rect 13589 275807 13623 275835
rect 13651 275807 13699 275835
rect 13389 275773 13699 275807
rect 13389 275745 13437 275773
rect 13465 275745 13499 275773
rect 13527 275745 13561 275773
rect 13589 275745 13623 275773
rect 13651 275745 13699 275773
rect 13389 266959 13699 275745
rect 13389 266931 13437 266959
rect 13465 266931 13499 266959
rect 13527 266931 13561 266959
rect 13589 266931 13623 266959
rect 13651 266931 13699 266959
rect 13389 266897 13699 266931
rect 13389 266869 13437 266897
rect 13465 266869 13499 266897
rect 13527 266869 13561 266897
rect 13589 266869 13623 266897
rect 13651 266869 13699 266897
rect 13389 266835 13699 266869
rect 13389 266807 13437 266835
rect 13465 266807 13499 266835
rect 13527 266807 13561 266835
rect 13589 266807 13623 266835
rect 13651 266807 13699 266835
rect 13389 266773 13699 266807
rect 13389 266745 13437 266773
rect 13465 266745 13499 266773
rect 13527 266745 13561 266773
rect 13589 266745 13623 266773
rect 13651 266745 13699 266773
rect 13389 257959 13699 266745
rect 13389 257931 13437 257959
rect 13465 257931 13499 257959
rect 13527 257931 13561 257959
rect 13589 257931 13623 257959
rect 13651 257931 13699 257959
rect 13389 257897 13699 257931
rect 13389 257869 13437 257897
rect 13465 257869 13499 257897
rect 13527 257869 13561 257897
rect 13589 257869 13623 257897
rect 13651 257869 13699 257897
rect 13389 257835 13699 257869
rect 13389 257807 13437 257835
rect 13465 257807 13499 257835
rect 13527 257807 13561 257835
rect 13589 257807 13623 257835
rect 13651 257807 13699 257835
rect 13389 257773 13699 257807
rect 13389 257745 13437 257773
rect 13465 257745 13499 257773
rect 13527 257745 13561 257773
rect 13589 257745 13623 257773
rect 13651 257745 13699 257773
rect 13389 248959 13699 257745
rect 20529 299190 20839 299718
rect 20529 299162 20577 299190
rect 20605 299162 20639 299190
rect 20667 299162 20701 299190
rect 20729 299162 20763 299190
rect 20791 299162 20839 299190
rect 20529 299128 20839 299162
rect 20529 299100 20577 299128
rect 20605 299100 20639 299128
rect 20667 299100 20701 299128
rect 20729 299100 20763 299128
rect 20791 299100 20839 299128
rect 20529 299066 20839 299100
rect 20529 299038 20577 299066
rect 20605 299038 20639 299066
rect 20667 299038 20701 299066
rect 20729 299038 20763 299066
rect 20791 299038 20839 299066
rect 20529 299004 20839 299038
rect 20529 298976 20577 299004
rect 20605 298976 20639 299004
rect 20667 298976 20701 299004
rect 20729 298976 20763 299004
rect 20791 298976 20839 299004
rect 20529 290959 20839 298976
rect 20529 290931 20577 290959
rect 20605 290931 20639 290959
rect 20667 290931 20701 290959
rect 20729 290931 20763 290959
rect 20791 290931 20839 290959
rect 20529 290897 20839 290931
rect 20529 290869 20577 290897
rect 20605 290869 20639 290897
rect 20667 290869 20701 290897
rect 20729 290869 20763 290897
rect 20791 290869 20839 290897
rect 20529 290835 20839 290869
rect 20529 290807 20577 290835
rect 20605 290807 20639 290835
rect 20667 290807 20701 290835
rect 20729 290807 20763 290835
rect 20791 290807 20839 290835
rect 20529 290773 20839 290807
rect 20529 290745 20577 290773
rect 20605 290745 20639 290773
rect 20667 290745 20701 290773
rect 20729 290745 20763 290773
rect 20791 290745 20839 290773
rect 20529 281959 20839 290745
rect 20529 281931 20577 281959
rect 20605 281931 20639 281959
rect 20667 281931 20701 281959
rect 20729 281931 20763 281959
rect 20791 281931 20839 281959
rect 20529 281897 20839 281931
rect 20529 281869 20577 281897
rect 20605 281869 20639 281897
rect 20667 281869 20701 281897
rect 20729 281869 20763 281897
rect 20791 281869 20839 281897
rect 20529 281835 20839 281869
rect 20529 281807 20577 281835
rect 20605 281807 20639 281835
rect 20667 281807 20701 281835
rect 20729 281807 20763 281835
rect 20791 281807 20839 281835
rect 20529 281773 20839 281807
rect 20529 281745 20577 281773
rect 20605 281745 20639 281773
rect 20667 281745 20701 281773
rect 20729 281745 20763 281773
rect 20791 281745 20839 281773
rect 20529 272959 20839 281745
rect 20529 272931 20577 272959
rect 20605 272931 20639 272959
rect 20667 272931 20701 272959
rect 20729 272931 20763 272959
rect 20791 272931 20839 272959
rect 20529 272897 20839 272931
rect 20529 272869 20577 272897
rect 20605 272869 20639 272897
rect 20667 272869 20701 272897
rect 20729 272869 20763 272897
rect 20791 272869 20839 272897
rect 20529 272835 20839 272869
rect 20529 272807 20577 272835
rect 20605 272807 20639 272835
rect 20667 272807 20701 272835
rect 20729 272807 20763 272835
rect 20791 272807 20839 272835
rect 20529 272773 20839 272807
rect 20529 272745 20577 272773
rect 20605 272745 20639 272773
rect 20667 272745 20701 272773
rect 20729 272745 20763 272773
rect 20791 272745 20839 272773
rect 20529 263959 20839 272745
rect 20529 263931 20577 263959
rect 20605 263931 20639 263959
rect 20667 263931 20701 263959
rect 20729 263931 20763 263959
rect 20791 263931 20839 263959
rect 20529 263897 20839 263931
rect 20529 263869 20577 263897
rect 20605 263869 20639 263897
rect 20667 263869 20701 263897
rect 20729 263869 20763 263897
rect 20791 263869 20839 263897
rect 20529 263835 20839 263869
rect 20529 263807 20577 263835
rect 20605 263807 20639 263835
rect 20667 263807 20701 263835
rect 20729 263807 20763 263835
rect 20791 263807 20839 263835
rect 20529 263773 20839 263807
rect 20529 263745 20577 263773
rect 20605 263745 20639 263773
rect 20667 263745 20701 263773
rect 20729 263745 20763 263773
rect 20791 263745 20839 263773
rect 15190 255402 15218 255407
rect 15190 253666 15218 255374
rect 15190 253633 15218 253638
rect 20529 254959 20839 263745
rect 20529 254931 20577 254959
rect 20605 254931 20639 254959
rect 20667 254931 20701 254959
rect 20729 254931 20763 254959
rect 20791 254931 20839 254959
rect 20529 254897 20839 254931
rect 20529 254869 20577 254897
rect 20605 254869 20639 254897
rect 20667 254869 20701 254897
rect 20729 254869 20763 254897
rect 20791 254869 20839 254897
rect 20529 254835 20839 254869
rect 20529 254807 20577 254835
rect 20605 254807 20639 254835
rect 20667 254807 20701 254835
rect 20729 254807 20763 254835
rect 20791 254807 20839 254835
rect 20529 254773 20839 254807
rect 20529 254745 20577 254773
rect 20605 254745 20639 254773
rect 20667 254745 20701 254773
rect 20729 254745 20763 254773
rect 20791 254745 20839 254773
rect 13389 248931 13437 248959
rect 13465 248931 13499 248959
rect 13527 248931 13561 248959
rect 13589 248931 13623 248959
rect 13651 248931 13699 248959
rect 13389 248897 13699 248931
rect 13389 248869 13437 248897
rect 13465 248869 13499 248897
rect 13527 248869 13561 248897
rect 13589 248869 13623 248897
rect 13651 248869 13699 248897
rect 13389 248835 13699 248869
rect 13389 248807 13437 248835
rect 13465 248807 13499 248835
rect 13527 248807 13561 248835
rect 13589 248807 13623 248835
rect 13651 248807 13699 248835
rect 13389 248773 13699 248807
rect 13389 248745 13437 248773
rect 13465 248745 13499 248773
rect 13527 248745 13561 248773
rect 13589 248745 13623 248773
rect 13651 248745 13699 248773
rect 13389 239959 13699 248745
rect 17224 245959 17384 245976
rect 17224 245931 17259 245959
rect 17287 245931 17321 245959
rect 17349 245931 17384 245959
rect 17224 245897 17384 245931
rect 17224 245869 17259 245897
rect 17287 245869 17321 245897
rect 17349 245869 17384 245897
rect 17224 245835 17384 245869
rect 17224 245807 17259 245835
rect 17287 245807 17321 245835
rect 17349 245807 17384 245835
rect 17224 245773 17384 245807
rect 17224 245745 17259 245773
rect 17287 245745 17321 245773
rect 17349 245745 17384 245773
rect 17224 245728 17384 245745
rect 20529 245959 20839 254745
rect 20529 245931 20577 245959
rect 20605 245931 20639 245959
rect 20667 245931 20701 245959
rect 20729 245931 20763 245959
rect 20791 245931 20839 245959
rect 20529 245897 20839 245931
rect 20529 245869 20577 245897
rect 20605 245869 20639 245897
rect 20667 245869 20701 245897
rect 20729 245869 20763 245897
rect 20791 245869 20839 245897
rect 20529 245835 20839 245869
rect 20529 245807 20577 245835
rect 20605 245807 20639 245835
rect 20667 245807 20701 245835
rect 20729 245807 20763 245835
rect 20791 245807 20839 245835
rect 20529 245773 20839 245807
rect 20529 245745 20577 245773
rect 20605 245745 20639 245773
rect 20667 245745 20701 245773
rect 20729 245745 20763 245773
rect 20791 245745 20839 245773
rect 13389 239931 13437 239959
rect 13465 239931 13499 239959
rect 13527 239931 13561 239959
rect 13589 239931 13623 239959
rect 13651 239931 13699 239959
rect 13389 239897 13699 239931
rect 13389 239869 13437 239897
rect 13465 239869 13499 239897
rect 13527 239869 13561 239897
rect 13589 239869 13623 239897
rect 13651 239869 13699 239897
rect 13389 239835 13699 239869
rect 13389 239807 13437 239835
rect 13465 239807 13499 239835
rect 13527 239807 13561 239835
rect 13589 239807 13623 239835
rect 13651 239807 13699 239835
rect 13389 239773 13699 239807
rect 13389 239745 13437 239773
rect 13465 239745 13499 239773
rect 13527 239745 13561 239773
rect 13589 239745 13623 239773
rect 13651 239745 13699 239773
rect 13389 230959 13699 239745
rect 17224 236959 17384 236976
rect 17224 236931 17259 236959
rect 17287 236931 17321 236959
rect 17349 236931 17384 236959
rect 17224 236897 17384 236931
rect 17224 236869 17259 236897
rect 17287 236869 17321 236897
rect 17349 236869 17384 236897
rect 17224 236835 17384 236869
rect 17224 236807 17259 236835
rect 17287 236807 17321 236835
rect 17349 236807 17384 236835
rect 17224 236773 17384 236807
rect 17224 236745 17259 236773
rect 17287 236745 17321 236773
rect 17349 236745 17384 236773
rect 17224 236728 17384 236745
rect 20529 236959 20839 245745
rect 20529 236931 20577 236959
rect 20605 236931 20639 236959
rect 20667 236931 20701 236959
rect 20729 236931 20763 236959
rect 20791 236931 20839 236959
rect 20529 236897 20839 236931
rect 20529 236869 20577 236897
rect 20605 236869 20639 236897
rect 20667 236869 20701 236897
rect 20729 236869 20763 236897
rect 20791 236869 20839 236897
rect 20529 236835 20839 236869
rect 20529 236807 20577 236835
rect 20605 236807 20639 236835
rect 20667 236807 20701 236835
rect 20729 236807 20763 236835
rect 20791 236807 20839 236835
rect 20529 236773 20839 236807
rect 20529 236745 20577 236773
rect 20605 236745 20639 236773
rect 20667 236745 20701 236773
rect 20729 236745 20763 236773
rect 20791 236745 20839 236773
rect 13389 230931 13437 230959
rect 13465 230931 13499 230959
rect 13527 230931 13561 230959
rect 13589 230931 13623 230959
rect 13651 230931 13699 230959
rect 13389 230897 13699 230931
rect 13389 230869 13437 230897
rect 13465 230869 13499 230897
rect 13527 230869 13561 230897
rect 13589 230869 13623 230897
rect 13651 230869 13699 230897
rect 13389 230835 13699 230869
rect 13389 230807 13437 230835
rect 13465 230807 13499 230835
rect 13527 230807 13561 230835
rect 13589 230807 13623 230835
rect 13651 230807 13699 230835
rect 13389 230773 13699 230807
rect 13389 230745 13437 230773
rect 13465 230745 13499 230773
rect 13527 230745 13561 230773
rect 13589 230745 13623 230773
rect 13651 230745 13699 230773
rect 13389 221959 13699 230745
rect 17224 227959 17384 227976
rect 17224 227931 17259 227959
rect 17287 227931 17321 227959
rect 17349 227931 17384 227959
rect 17224 227897 17384 227931
rect 17224 227869 17259 227897
rect 17287 227869 17321 227897
rect 17349 227869 17384 227897
rect 17224 227835 17384 227869
rect 17224 227807 17259 227835
rect 17287 227807 17321 227835
rect 17349 227807 17384 227835
rect 17224 227773 17384 227807
rect 17224 227745 17259 227773
rect 17287 227745 17321 227773
rect 17349 227745 17384 227773
rect 17224 227728 17384 227745
rect 20529 227959 20839 236745
rect 20529 227931 20577 227959
rect 20605 227931 20639 227959
rect 20667 227931 20701 227959
rect 20729 227931 20763 227959
rect 20791 227931 20839 227959
rect 20529 227897 20839 227931
rect 20529 227869 20577 227897
rect 20605 227869 20639 227897
rect 20667 227869 20701 227897
rect 20729 227869 20763 227897
rect 20791 227869 20839 227897
rect 20529 227835 20839 227869
rect 20529 227807 20577 227835
rect 20605 227807 20639 227835
rect 20667 227807 20701 227835
rect 20729 227807 20763 227835
rect 20791 227807 20839 227835
rect 20529 227773 20839 227807
rect 20529 227745 20577 227773
rect 20605 227745 20639 227773
rect 20667 227745 20701 227773
rect 20729 227745 20763 227773
rect 20791 227745 20839 227773
rect 13389 221931 13437 221959
rect 13465 221931 13499 221959
rect 13527 221931 13561 221959
rect 13589 221931 13623 221959
rect 13651 221931 13699 221959
rect 13389 221897 13699 221931
rect 13389 221869 13437 221897
rect 13465 221869 13499 221897
rect 13527 221869 13561 221897
rect 13589 221869 13623 221897
rect 13651 221869 13699 221897
rect 13389 221835 13699 221869
rect 13389 221807 13437 221835
rect 13465 221807 13499 221835
rect 13527 221807 13561 221835
rect 13589 221807 13623 221835
rect 13651 221807 13699 221835
rect 13389 221773 13699 221807
rect 13389 221745 13437 221773
rect 13465 221745 13499 221773
rect 13527 221745 13561 221773
rect 13589 221745 13623 221773
rect 13651 221745 13699 221773
rect 13389 212959 13699 221745
rect 17224 218959 17384 218976
rect 17224 218931 17259 218959
rect 17287 218931 17321 218959
rect 17349 218931 17384 218959
rect 17224 218897 17384 218931
rect 17224 218869 17259 218897
rect 17287 218869 17321 218897
rect 17349 218869 17384 218897
rect 17224 218835 17384 218869
rect 17224 218807 17259 218835
rect 17287 218807 17321 218835
rect 17349 218807 17384 218835
rect 17224 218773 17384 218807
rect 17224 218745 17259 218773
rect 17287 218745 17321 218773
rect 17349 218745 17384 218773
rect 17224 218728 17384 218745
rect 20529 218959 20839 227745
rect 20529 218931 20577 218959
rect 20605 218931 20639 218959
rect 20667 218931 20701 218959
rect 20729 218931 20763 218959
rect 20791 218931 20839 218959
rect 20529 218897 20839 218931
rect 20529 218869 20577 218897
rect 20605 218869 20639 218897
rect 20667 218869 20701 218897
rect 20729 218869 20763 218897
rect 20791 218869 20839 218897
rect 20529 218835 20839 218869
rect 20529 218807 20577 218835
rect 20605 218807 20639 218835
rect 20667 218807 20701 218835
rect 20729 218807 20763 218835
rect 20791 218807 20839 218835
rect 20529 218773 20839 218807
rect 20529 218745 20577 218773
rect 20605 218745 20639 218773
rect 20667 218745 20701 218773
rect 20729 218745 20763 218773
rect 20791 218745 20839 218773
rect 13389 212931 13437 212959
rect 13465 212931 13499 212959
rect 13527 212931 13561 212959
rect 13589 212931 13623 212959
rect 13651 212931 13699 212959
rect 13389 212897 13699 212931
rect 13389 212869 13437 212897
rect 13465 212869 13499 212897
rect 13527 212869 13561 212897
rect 13589 212869 13623 212897
rect 13651 212869 13699 212897
rect 13389 212835 13699 212869
rect 13389 212807 13437 212835
rect 13465 212807 13499 212835
rect 13527 212807 13561 212835
rect 13589 212807 13623 212835
rect 13651 212807 13699 212835
rect 13389 212773 13699 212807
rect 13389 212745 13437 212773
rect 13465 212745 13499 212773
rect 13527 212745 13561 212773
rect 13589 212745 13623 212773
rect 13651 212745 13699 212773
rect 13389 203959 13699 212745
rect 17224 209959 17384 209976
rect 17224 209931 17259 209959
rect 17287 209931 17321 209959
rect 17349 209931 17384 209959
rect 17224 209897 17384 209931
rect 17224 209869 17259 209897
rect 17287 209869 17321 209897
rect 17349 209869 17384 209897
rect 17224 209835 17384 209869
rect 17224 209807 17259 209835
rect 17287 209807 17321 209835
rect 17349 209807 17384 209835
rect 17224 209773 17384 209807
rect 17224 209745 17259 209773
rect 17287 209745 17321 209773
rect 17349 209745 17384 209773
rect 17224 209728 17384 209745
rect 20529 209959 20839 218745
rect 20529 209931 20577 209959
rect 20605 209931 20639 209959
rect 20667 209931 20701 209959
rect 20729 209931 20763 209959
rect 20791 209931 20839 209959
rect 20529 209897 20839 209931
rect 20529 209869 20577 209897
rect 20605 209869 20639 209897
rect 20667 209869 20701 209897
rect 20729 209869 20763 209897
rect 20791 209869 20839 209897
rect 20529 209835 20839 209869
rect 20529 209807 20577 209835
rect 20605 209807 20639 209835
rect 20667 209807 20701 209835
rect 20729 209807 20763 209835
rect 20791 209807 20839 209835
rect 20529 209773 20839 209807
rect 20529 209745 20577 209773
rect 20605 209745 20639 209773
rect 20667 209745 20701 209773
rect 20729 209745 20763 209773
rect 20791 209745 20839 209773
rect 13389 203931 13437 203959
rect 13465 203931 13499 203959
rect 13527 203931 13561 203959
rect 13589 203931 13623 203959
rect 13651 203931 13699 203959
rect 13389 203897 13699 203931
rect 13389 203869 13437 203897
rect 13465 203869 13499 203897
rect 13527 203869 13561 203897
rect 13589 203869 13623 203897
rect 13651 203869 13699 203897
rect 13389 203835 13699 203869
rect 13389 203807 13437 203835
rect 13465 203807 13499 203835
rect 13527 203807 13561 203835
rect 13589 203807 13623 203835
rect 13651 203807 13699 203835
rect 13389 203773 13699 203807
rect 13389 203745 13437 203773
rect 13465 203745 13499 203773
rect 13527 203745 13561 203773
rect 13589 203745 13623 203773
rect 13651 203745 13699 203773
rect 13389 194959 13699 203745
rect 17224 200959 17384 200976
rect 17224 200931 17259 200959
rect 17287 200931 17321 200959
rect 17349 200931 17384 200959
rect 17224 200897 17384 200931
rect 17224 200869 17259 200897
rect 17287 200869 17321 200897
rect 17349 200869 17384 200897
rect 17224 200835 17384 200869
rect 17224 200807 17259 200835
rect 17287 200807 17321 200835
rect 17349 200807 17384 200835
rect 17224 200773 17384 200807
rect 17224 200745 17259 200773
rect 17287 200745 17321 200773
rect 17349 200745 17384 200773
rect 17224 200728 17384 200745
rect 20529 200959 20839 209745
rect 20529 200931 20577 200959
rect 20605 200931 20639 200959
rect 20667 200931 20701 200959
rect 20729 200931 20763 200959
rect 20791 200931 20839 200959
rect 20529 200897 20839 200931
rect 20529 200869 20577 200897
rect 20605 200869 20639 200897
rect 20667 200869 20701 200897
rect 20729 200869 20763 200897
rect 20791 200869 20839 200897
rect 20529 200835 20839 200869
rect 20529 200807 20577 200835
rect 20605 200807 20639 200835
rect 20667 200807 20701 200835
rect 20729 200807 20763 200835
rect 20791 200807 20839 200835
rect 20529 200773 20839 200807
rect 20529 200745 20577 200773
rect 20605 200745 20639 200773
rect 20667 200745 20701 200773
rect 20729 200745 20763 200773
rect 20791 200745 20839 200773
rect 13389 194931 13437 194959
rect 13465 194931 13499 194959
rect 13527 194931 13561 194959
rect 13589 194931 13623 194959
rect 13651 194931 13699 194959
rect 13389 194897 13699 194931
rect 13389 194869 13437 194897
rect 13465 194869 13499 194897
rect 13527 194869 13561 194897
rect 13589 194869 13623 194897
rect 13651 194869 13699 194897
rect 13389 194835 13699 194869
rect 13389 194807 13437 194835
rect 13465 194807 13499 194835
rect 13527 194807 13561 194835
rect 13589 194807 13623 194835
rect 13651 194807 13699 194835
rect 13389 194773 13699 194807
rect 13389 194745 13437 194773
rect 13465 194745 13499 194773
rect 13527 194745 13561 194773
rect 13589 194745 13623 194773
rect 13651 194745 13699 194773
rect 13389 185959 13699 194745
rect 17224 191959 17384 191976
rect 17224 191931 17259 191959
rect 17287 191931 17321 191959
rect 17349 191931 17384 191959
rect 17224 191897 17384 191931
rect 17224 191869 17259 191897
rect 17287 191869 17321 191897
rect 17349 191869 17384 191897
rect 17224 191835 17384 191869
rect 17224 191807 17259 191835
rect 17287 191807 17321 191835
rect 17349 191807 17384 191835
rect 17224 191773 17384 191807
rect 17224 191745 17259 191773
rect 17287 191745 17321 191773
rect 17349 191745 17384 191773
rect 17224 191728 17384 191745
rect 20529 191959 20839 200745
rect 20529 191931 20577 191959
rect 20605 191931 20639 191959
rect 20667 191931 20701 191959
rect 20729 191931 20763 191959
rect 20791 191931 20839 191959
rect 20529 191897 20839 191931
rect 20529 191869 20577 191897
rect 20605 191869 20639 191897
rect 20667 191869 20701 191897
rect 20729 191869 20763 191897
rect 20791 191869 20839 191897
rect 20529 191835 20839 191869
rect 20529 191807 20577 191835
rect 20605 191807 20639 191835
rect 20667 191807 20701 191835
rect 20729 191807 20763 191835
rect 20791 191807 20839 191835
rect 20529 191773 20839 191807
rect 20529 191745 20577 191773
rect 20605 191745 20639 191773
rect 20667 191745 20701 191773
rect 20729 191745 20763 191773
rect 20791 191745 20839 191773
rect 13389 185931 13437 185959
rect 13465 185931 13499 185959
rect 13527 185931 13561 185959
rect 13589 185931 13623 185959
rect 13651 185931 13699 185959
rect 13389 185897 13699 185931
rect 13389 185869 13437 185897
rect 13465 185869 13499 185897
rect 13527 185869 13561 185897
rect 13589 185869 13623 185897
rect 13651 185869 13699 185897
rect 13389 185835 13699 185869
rect 13389 185807 13437 185835
rect 13465 185807 13499 185835
rect 13527 185807 13561 185835
rect 13589 185807 13623 185835
rect 13651 185807 13699 185835
rect 13389 185773 13699 185807
rect 13389 185745 13437 185773
rect 13465 185745 13499 185773
rect 13527 185745 13561 185773
rect 13589 185745 13623 185773
rect 13651 185745 13699 185773
rect 13389 176959 13699 185745
rect 17224 182959 17384 182976
rect 17224 182931 17259 182959
rect 17287 182931 17321 182959
rect 17349 182931 17384 182959
rect 17224 182897 17384 182931
rect 17224 182869 17259 182897
rect 17287 182869 17321 182897
rect 17349 182869 17384 182897
rect 17224 182835 17384 182869
rect 17224 182807 17259 182835
rect 17287 182807 17321 182835
rect 17349 182807 17384 182835
rect 17224 182773 17384 182807
rect 17224 182745 17259 182773
rect 17287 182745 17321 182773
rect 17349 182745 17384 182773
rect 17224 182728 17384 182745
rect 20529 182959 20839 191745
rect 20529 182931 20577 182959
rect 20605 182931 20639 182959
rect 20667 182931 20701 182959
rect 20729 182931 20763 182959
rect 20791 182931 20839 182959
rect 20529 182897 20839 182931
rect 20529 182869 20577 182897
rect 20605 182869 20639 182897
rect 20667 182869 20701 182897
rect 20729 182869 20763 182897
rect 20791 182869 20839 182897
rect 20529 182835 20839 182869
rect 20529 182807 20577 182835
rect 20605 182807 20639 182835
rect 20667 182807 20701 182835
rect 20729 182807 20763 182835
rect 20791 182807 20839 182835
rect 20529 182773 20839 182807
rect 20529 182745 20577 182773
rect 20605 182745 20639 182773
rect 20667 182745 20701 182773
rect 20729 182745 20763 182773
rect 20791 182745 20839 182773
rect 13389 176931 13437 176959
rect 13465 176931 13499 176959
rect 13527 176931 13561 176959
rect 13589 176931 13623 176959
rect 13651 176931 13699 176959
rect 13389 176897 13699 176931
rect 13389 176869 13437 176897
rect 13465 176869 13499 176897
rect 13527 176869 13561 176897
rect 13589 176869 13623 176897
rect 13651 176869 13699 176897
rect 13389 176835 13699 176869
rect 13389 176807 13437 176835
rect 13465 176807 13499 176835
rect 13527 176807 13561 176835
rect 13589 176807 13623 176835
rect 13651 176807 13699 176835
rect 13389 176773 13699 176807
rect 13389 176745 13437 176773
rect 13465 176745 13499 176773
rect 13527 176745 13561 176773
rect 13589 176745 13623 176773
rect 13651 176745 13699 176773
rect 13389 167959 13699 176745
rect 17224 173959 17384 173976
rect 17224 173931 17259 173959
rect 17287 173931 17321 173959
rect 17349 173931 17384 173959
rect 17224 173897 17384 173931
rect 17224 173869 17259 173897
rect 17287 173869 17321 173897
rect 17349 173869 17384 173897
rect 17224 173835 17384 173869
rect 17224 173807 17259 173835
rect 17287 173807 17321 173835
rect 17349 173807 17384 173835
rect 17224 173773 17384 173807
rect 17224 173745 17259 173773
rect 17287 173745 17321 173773
rect 17349 173745 17384 173773
rect 17224 173728 17384 173745
rect 20529 173959 20839 182745
rect 20529 173931 20577 173959
rect 20605 173931 20639 173959
rect 20667 173931 20701 173959
rect 20729 173931 20763 173959
rect 20791 173931 20839 173959
rect 20529 173897 20839 173931
rect 20529 173869 20577 173897
rect 20605 173869 20639 173897
rect 20667 173869 20701 173897
rect 20729 173869 20763 173897
rect 20791 173869 20839 173897
rect 20529 173835 20839 173869
rect 20529 173807 20577 173835
rect 20605 173807 20639 173835
rect 20667 173807 20701 173835
rect 20729 173807 20763 173835
rect 20791 173807 20839 173835
rect 20529 173773 20839 173807
rect 20529 173745 20577 173773
rect 20605 173745 20639 173773
rect 20667 173745 20701 173773
rect 20729 173745 20763 173773
rect 20791 173745 20839 173773
rect 13389 167931 13437 167959
rect 13465 167931 13499 167959
rect 13527 167931 13561 167959
rect 13589 167931 13623 167959
rect 13651 167931 13699 167959
rect 13389 167897 13699 167931
rect 13389 167869 13437 167897
rect 13465 167869 13499 167897
rect 13527 167869 13561 167897
rect 13589 167869 13623 167897
rect 13651 167869 13699 167897
rect 13389 167835 13699 167869
rect 13389 167807 13437 167835
rect 13465 167807 13499 167835
rect 13527 167807 13561 167835
rect 13589 167807 13623 167835
rect 13651 167807 13699 167835
rect 13389 167773 13699 167807
rect 13389 167745 13437 167773
rect 13465 167745 13499 167773
rect 13527 167745 13561 167773
rect 13589 167745 13623 167773
rect 13651 167745 13699 167773
rect 13389 158959 13699 167745
rect 17224 164959 17384 164976
rect 17224 164931 17259 164959
rect 17287 164931 17321 164959
rect 17349 164931 17384 164959
rect 17224 164897 17384 164931
rect 17224 164869 17259 164897
rect 17287 164869 17321 164897
rect 17349 164869 17384 164897
rect 17224 164835 17384 164869
rect 17224 164807 17259 164835
rect 17287 164807 17321 164835
rect 17349 164807 17384 164835
rect 17224 164773 17384 164807
rect 17224 164745 17259 164773
rect 17287 164745 17321 164773
rect 17349 164745 17384 164773
rect 17224 164728 17384 164745
rect 20529 164959 20839 173745
rect 20529 164931 20577 164959
rect 20605 164931 20639 164959
rect 20667 164931 20701 164959
rect 20729 164931 20763 164959
rect 20791 164931 20839 164959
rect 20529 164897 20839 164931
rect 20529 164869 20577 164897
rect 20605 164869 20639 164897
rect 20667 164869 20701 164897
rect 20729 164869 20763 164897
rect 20791 164869 20839 164897
rect 20529 164835 20839 164869
rect 20529 164807 20577 164835
rect 20605 164807 20639 164835
rect 20667 164807 20701 164835
rect 20729 164807 20763 164835
rect 20791 164807 20839 164835
rect 20529 164773 20839 164807
rect 20529 164745 20577 164773
rect 20605 164745 20639 164773
rect 20667 164745 20701 164773
rect 20729 164745 20763 164773
rect 20791 164745 20839 164773
rect 13389 158931 13437 158959
rect 13465 158931 13499 158959
rect 13527 158931 13561 158959
rect 13589 158931 13623 158959
rect 13651 158931 13699 158959
rect 13389 158897 13699 158931
rect 13389 158869 13437 158897
rect 13465 158869 13499 158897
rect 13527 158869 13561 158897
rect 13589 158869 13623 158897
rect 13651 158869 13699 158897
rect 13389 158835 13699 158869
rect 13389 158807 13437 158835
rect 13465 158807 13499 158835
rect 13527 158807 13561 158835
rect 13589 158807 13623 158835
rect 13651 158807 13699 158835
rect 13389 158773 13699 158807
rect 13389 158745 13437 158773
rect 13465 158745 13499 158773
rect 13527 158745 13561 158773
rect 13589 158745 13623 158773
rect 13651 158745 13699 158773
rect 13389 149959 13699 158745
rect 17224 155959 17384 155976
rect 17224 155931 17259 155959
rect 17287 155931 17321 155959
rect 17349 155931 17384 155959
rect 17224 155897 17384 155931
rect 17224 155869 17259 155897
rect 17287 155869 17321 155897
rect 17349 155869 17384 155897
rect 17224 155835 17384 155869
rect 17224 155807 17259 155835
rect 17287 155807 17321 155835
rect 17349 155807 17384 155835
rect 17224 155773 17384 155807
rect 17224 155745 17259 155773
rect 17287 155745 17321 155773
rect 17349 155745 17384 155773
rect 17224 155728 17384 155745
rect 20529 155959 20839 164745
rect 20529 155931 20577 155959
rect 20605 155931 20639 155959
rect 20667 155931 20701 155959
rect 20729 155931 20763 155959
rect 20791 155931 20839 155959
rect 20529 155897 20839 155931
rect 20529 155869 20577 155897
rect 20605 155869 20639 155897
rect 20667 155869 20701 155897
rect 20729 155869 20763 155897
rect 20791 155869 20839 155897
rect 20529 155835 20839 155869
rect 20529 155807 20577 155835
rect 20605 155807 20639 155835
rect 20667 155807 20701 155835
rect 20729 155807 20763 155835
rect 20791 155807 20839 155835
rect 20529 155773 20839 155807
rect 20529 155745 20577 155773
rect 20605 155745 20639 155773
rect 20667 155745 20701 155773
rect 20729 155745 20763 155773
rect 20791 155745 20839 155773
rect 13389 149931 13437 149959
rect 13465 149931 13499 149959
rect 13527 149931 13561 149959
rect 13589 149931 13623 149959
rect 13651 149931 13699 149959
rect 13389 149897 13699 149931
rect 13389 149869 13437 149897
rect 13465 149869 13499 149897
rect 13527 149869 13561 149897
rect 13589 149869 13623 149897
rect 13651 149869 13699 149897
rect 13389 149835 13699 149869
rect 13389 149807 13437 149835
rect 13465 149807 13499 149835
rect 13527 149807 13561 149835
rect 13589 149807 13623 149835
rect 13651 149807 13699 149835
rect 13389 149773 13699 149807
rect 13389 149745 13437 149773
rect 13465 149745 13499 149773
rect 13527 149745 13561 149773
rect 13589 149745 13623 149773
rect 13651 149745 13699 149773
rect 13389 140959 13699 149745
rect 17224 146959 17384 146976
rect 17224 146931 17259 146959
rect 17287 146931 17321 146959
rect 17349 146931 17384 146959
rect 17224 146897 17384 146931
rect 17224 146869 17259 146897
rect 17287 146869 17321 146897
rect 17349 146869 17384 146897
rect 17224 146835 17384 146869
rect 17224 146807 17259 146835
rect 17287 146807 17321 146835
rect 17349 146807 17384 146835
rect 17224 146773 17384 146807
rect 17224 146745 17259 146773
rect 17287 146745 17321 146773
rect 17349 146745 17384 146773
rect 17224 146728 17384 146745
rect 20529 146959 20839 155745
rect 20529 146931 20577 146959
rect 20605 146931 20639 146959
rect 20667 146931 20701 146959
rect 20729 146931 20763 146959
rect 20791 146931 20839 146959
rect 20529 146897 20839 146931
rect 20529 146869 20577 146897
rect 20605 146869 20639 146897
rect 20667 146869 20701 146897
rect 20729 146869 20763 146897
rect 20791 146869 20839 146897
rect 20529 146835 20839 146869
rect 20529 146807 20577 146835
rect 20605 146807 20639 146835
rect 20667 146807 20701 146835
rect 20729 146807 20763 146835
rect 20791 146807 20839 146835
rect 20529 146773 20839 146807
rect 20529 146745 20577 146773
rect 20605 146745 20639 146773
rect 20667 146745 20701 146773
rect 20729 146745 20763 146773
rect 20791 146745 20839 146773
rect 13389 140931 13437 140959
rect 13465 140931 13499 140959
rect 13527 140931 13561 140959
rect 13589 140931 13623 140959
rect 13651 140931 13699 140959
rect 13389 140897 13699 140931
rect 13389 140869 13437 140897
rect 13465 140869 13499 140897
rect 13527 140869 13561 140897
rect 13589 140869 13623 140897
rect 13651 140869 13699 140897
rect 13389 140835 13699 140869
rect 13389 140807 13437 140835
rect 13465 140807 13499 140835
rect 13527 140807 13561 140835
rect 13589 140807 13623 140835
rect 13651 140807 13699 140835
rect 13389 140773 13699 140807
rect 13389 140745 13437 140773
rect 13465 140745 13499 140773
rect 13527 140745 13561 140773
rect 13589 140745 13623 140773
rect 13651 140745 13699 140773
rect 13389 131959 13699 140745
rect 17224 137959 17384 137976
rect 17224 137931 17259 137959
rect 17287 137931 17321 137959
rect 17349 137931 17384 137959
rect 17224 137897 17384 137931
rect 17224 137869 17259 137897
rect 17287 137869 17321 137897
rect 17349 137869 17384 137897
rect 17224 137835 17384 137869
rect 17224 137807 17259 137835
rect 17287 137807 17321 137835
rect 17349 137807 17384 137835
rect 17224 137773 17384 137807
rect 17224 137745 17259 137773
rect 17287 137745 17321 137773
rect 17349 137745 17384 137773
rect 17224 137728 17384 137745
rect 20529 137959 20839 146745
rect 20529 137931 20577 137959
rect 20605 137931 20639 137959
rect 20667 137931 20701 137959
rect 20729 137931 20763 137959
rect 20791 137931 20839 137959
rect 20529 137897 20839 137931
rect 20529 137869 20577 137897
rect 20605 137869 20639 137897
rect 20667 137869 20701 137897
rect 20729 137869 20763 137897
rect 20791 137869 20839 137897
rect 20529 137835 20839 137869
rect 20529 137807 20577 137835
rect 20605 137807 20639 137835
rect 20667 137807 20701 137835
rect 20729 137807 20763 137835
rect 20791 137807 20839 137835
rect 20529 137773 20839 137807
rect 20529 137745 20577 137773
rect 20605 137745 20639 137773
rect 20667 137745 20701 137773
rect 20729 137745 20763 137773
rect 20791 137745 20839 137773
rect 13389 131931 13437 131959
rect 13465 131931 13499 131959
rect 13527 131931 13561 131959
rect 13589 131931 13623 131959
rect 13651 131931 13699 131959
rect 13389 131897 13699 131931
rect 13389 131869 13437 131897
rect 13465 131869 13499 131897
rect 13527 131869 13561 131897
rect 13589 131869 13623 131897
rect 13651 131869 13699 131897
rect 13389 131835 13699 131869
rect 13389 131807 13437 131835
rect 13465 131807 13499 131835
rect 13527 131807 13561 131835
rect 13589 131807 13623 131835
rect 13651 131807 13699 131835
rect 13389 131773 13699 131807
rect 13389 131745 13437 131773
rect 13465 131745 13499 131773
rect 13527 131745 13561 131773
rect 13589 131745 13623 131773
rect 13651 131745 13699 131773
rect 13389 122959 13699 131745
rect 17224 128959 17384 128976
rect 17224 128931 17259 128959
rect 17287 128931 17321 128959
rect 17349 128931 17384 128959
rect 17224 128897 17384 128931
rect 17224 128869 17259 128897
rect 17287 128869 17321 128897
rect 17349 128869 17384 128897
rect 17224 128835 17384 128869
rect 17224 128807 17259 128835
rect 17287 128807 17321 128835
rect 17349 128807 17384 128835
rect 17224 128773 17384 128807
rect 17224 128745 17259 128773
rect 17287 128745 17321 128773
rect 17349 128745 17384 128773
rect 17224 128728 17384 128745
rect 20529 128959 20839 137745
rect 20529 128931 20577 128959
rect 20605 128931 20639 128959
rect 20667 128931 20701 128959
rect 20729 128931 20763 128959
rect 20791 128931 20839 128959
rect 20529 128897 20839 128931
rect 20529 128869 20577 128897
rect 20605 128869 20639 128897
rect 20667 128869 20701 128897
rect 20729 128869 20763 128897
rect 20791 128869 20839 128897
rect 20529 128835 20839 128869
rect 20529 128807 20577 128835
rect 20605 128807 20639 128835
rect 20667 128807 20701 128835
rect 20729 128807 20763 128835
rect 20791 128807 20839 128835
rect 20529 128773 20839 128807
rect 20529 128745 20577 128773
rect 20605 128745 20639 128773
rect 20667 128745 20701 128773
rect 20729 128745 20763 128773
rect 20791 128745 20839 128773
rect 13389 122931 13437 122959
rect 13465 122931 13499 122959
rect 13527 122931 13561 122959
rect 13589 122931 13623 122959
rect 13651 122931 13699 122959
rect 13389 122897 13699 122931
rect 13389 122869 13437 122897
rect 13465 122869 13499 122897
rect 13527 122869 13561 122897
rect 13589 122869 13623 122897
rect 13651 122869 13699 122897
rect 13389 122835 13699 122869
rect 13389 122807 13437 122835
rect 13465 122807 13499 122835
rect 13527 122807 13561 122835
rect 13589 122807 13623 122835
rect 13651 122807 13699 122835
rect 13389 122773 13699 122807
rect 13389 122745 13437 122773
rect 13465 122745 13499 122773
rect 13527 122745 13561 122773
rect 13589 122745 13623 122773
rect 13651 122745 13699 122773
rect 13389 113959 13699 122745
rect 17224 119959 17384 119976
rect 17224 119931 17259 119959
rect 17287 119931 17321 119959
rect 17349 119931 17384 119959
rect 17224 119897 17384 119931
rect 17224 119869 17259 119897
rect 17287 119869 17321 119897
rect 17349 119869 17384 119897
rect 17224 119835 17384 119869
rect 17224 119807 17259 119835
rect 17287 119807 17321 119835
rect 17349 119807 17384 119835
rect 17224 119773 17384 119807
rect 17224 119745 17259 119773
rect 17287 119745 17321 119773
rect 17349 119745 17384 119773
rect 17224 119728 17384 119745
rect 20529 119959 20839 128745
rect 20529 119931 20577 119959
rect 20605 119931 20639 119959
rect 20667 119931 20701 119959
rect 20729 119931 20763 119959
rect 20791 119931 20839 119959
rect 20529 119897 20839 119931
rect 20529 119869 20577 119897
rect 20605 119869 20639 119897
rect 20667 119869 20701 119897
rect 20729 119869 20763 119897
rect 20791 119869 20839 119897
rect 20529 119835 20839 119869
rect 20529 119807 20577 119835
rect 20605 119807 20639 119835
rect 20667 119807 20701 119835
rect 20729 119807 20763 119835
rect 20791 119807 20839 119835
rect 20529 119773 20839 119807
rect 20529 119745 20577 119773
rect 20605 119745 20639 119773
rect 20667 119745 20701 119773
rect 20729 119745 20763 119773
rect 20791 119745 20839 119773
rect 13389 113931 13437 113959
rect 13465 113931 13499 113959
rect 13527 113931 13561 113959
rect 13589 113931 13623 113959
rect 13651 113931 13699 113959
rect 13389 113897 13699 113931
rect 13389 113869 13437 113897
rect 13465 113869 13499 113897
rect 13527 113869 13561 113897
rect 13589 113869 13623 113897
rect 13651 113869 13699 113897
rect 13389 113835 13699 113869
rect 13389 113807 13437 113835
rect 13465 113807 13499 113835
rect 13527 113807 13561 113835
rect 13589 113807 13623 113835
rect 13651 113807 13699 113835
rect 13389 113773 13699 113807
rect 13389 113745 13437 113773
rect 13465 113745 13499 113773
rect 13527 113745 13561 113773
rect 13589 113745 13623 113773
rect 13651 113745 13699 113773
rect 13389 104959 13699 113745
rect 17224 110959 17384 110976
rect 17224 110931 17259 110959
rect 17287 110931 17321 110959
rect 17349 110931 17384 110959
rect 17224 110897 17384 110931
rect 17224 110869 17259 110897
rect 17287 110869 17321 110897
rect 17349 110869 17384 110897
rect 17224 110835 17384 110869
rect 17224 110807 17259 110835
rect 17287 110807 17321 110835
rect 17349 110807 17384 110835
rect 17224 110773 17384 110807
rect 17224 110745 17259 110773
rect 17287 110745 17321 110773
rect 17349 110745 17384 110773
rect 17224 110728 17384 110745
rect 20529 110959 20839 119745
rect 20529 110931 20577 110959
rect 20605 110931 20639 110959
rect 20667 110931 20701 110959
rect 20729 110931 20763 110959
rect 20791 110931 20839 110959
rect 20529 110897 20839 110931
rect 20529 110869 20577 110897
rect 20605 110869 20639 110897
rect 20667 110869 20701 110897
rect 20729 110869 20763 110897
rect 20791 110869 20839 110897
rect 20529 110835 20839 110869
rect 20529 110807 20577 110835
rect 20605 110807 20639 110835
rect 20667 110807 20701 110835
rect 20729 110807 20763 110835
rect 20791 110807 20839 110835
rect 20529 110773 20839 110807
rect 20529 110745 20577 110773
rect 20605 110745 20639 110773
rect 20667 110745 20701 110773
rect 20729 110745 20763 110773
rect 20791 110745 20839 110773
rect 13389 104931 13437 104959
rect 13465 104931 13499 104959
rect 13527 104931 13561 104959
rect 13589 104931 13623 104959
rect 13651 104931 13699 104959
rect 13389 104897 13699 104931
rect 13389 104869 13437 104897
rect 13465 104869 13499 104897
rect 13527 104869 13561 104897
rect 13589 104869 13623 104897
rect 13651 104869 13699 104897
rect 13389 104835 13699 104869
rect 13389 104807 13437 104835
rect 13465 104807 13499 104835
rect 13527 104807 13561 104835
rect 13589 104807 13623 104835
rect 13651 104807 13699 104835
rect 13389 104773 13699 104807
rect 13389 104745 13437 104773
rect 13465 104745 13499 104773
rect 13527 104745 13561 104773
rect 13589 104745 13623 104773
rect 13651 104745 13699 104773
rect 13389 95959 13699 104745
rect 17224 101959 17384 101976
rect 17224 101931 17259 101959
rect 17287 101931 17321 101959
rect 17349 101931 17384 101959
rect 17224 101897 17384 101931
rect 17224 101869 17259 101897
rect 17287 101869 17321 101897
rect 17349 101869 17384 101897
rect 17224 101835 17384 101869
rect 17224 101807 17259 101835
rect 17287 101807 17321 101835
rect 17349 101807 17384 101835
rect 17224 101773 17384 101807
rect 17224 101745 17259 101773
rect 17287 101745 17321 101773
rect 17349 101745 17384 101773
rect 17224 101728 17384 101745
rect 20529 101959 20839 110745
rect 20529 101931 20577 101959
rect 20605 101931 20639 101959
rect 20667 101931 20701 101959
rect 20729 101931 20763 101959
rect 20791 101931 20839 101959
rect 20529 101897 20839 101931
rect 20529 101869 20577 101897
rect 20605 101869 20639 101897
rect 20667 101869 20701 101897
rect 20729 101869 20763 101897
rect 20791 101869 20839 101897
rect 20529 101835 20839 101869
rect 20529 101807 20577 101835
rect 20605 101807 20639 101835
rect 20667 101807 20701 101835
rect 20729 101807 20763 101835
rect 20791 101807 20839 101835
rect 20529 101773 20839 101807
rect 20529 101745 20577 101773
rect 20605 101745 20639 101773
rect 20667 101745 20701 101773
rect 20729 101745 20763 101773
rect 20791 101745 20839 101773
rect 13389 95931 13437 95959
rect 13465 95931 13499 95959
rect 13527 95931 13561 95959
rect 13589 95931 13623 95959
rect 13651 95931 13699 95959
rect 13389 95897 13699 95931
rect 13389 95869 13437 95897
rect 13465 95869 13499 95897
rect 13527 95869 13561 95897
rect 13589 95869 13623 95897
rect 13651 95869 13699 95897
rect 13389 95835 13699 95869
rect 13389 95807 13437 95835
rect 13465 95807 13499 95835
rect 13527 95807 13561 95835
rect 13589 95807 13623 95835
rect 13651 95807 13699 95835
rect 13389 95773 13699 95807
rect 13389 95745 13437 95773
rect 13465 95745 13499 95773
rect 13527 95745 13561 95773
rect 13589 95745 13623 95773
rect 13651 95745 13699 95773
rect 13389 86959 13699 95745
rect 17224 92959 17384 92976
rect 17224 92931 17259 92959
rect 17287 92931 17321 92959
rect 17349 92931 17384 92959
rect 17224 92897 17384 92931
rect 17224 92869 17259 92897
rect 17287 92869 17321 92897
rect 17349 92869 17384 92897
rect 17224 92835 17384 92869
rect 17224 92807 17259 92835
rect 17287 92807 17321 92835
rect 17349 92807 17384 92835
rect 17224 92773 17384 92807
rect 17224 92745 17259 92773
rect 17287 92745 17321 92773
rect 17349 92745 17384 92773
rect 17224 92728 17384 92745
rect 20529 92959 20839 101745
rect 20529 92931 20577 92959
rect 20605 92931 20639 92959
rect 20667 92931 20701 92959
rect 20729 92931 20763 92959
rect 20791 92931 20839 92959
rect 20529 92897 20839 92931
rect 20529 92869 20577 92897
rect 20605 92869 20639 92897
rect 20667 92869 20701 92897
rect 20729 92869 20763 92897
rect 20791 92869 20839 92897
rect 20529 92835 20839 92869
rect 20529 92807 20577 92835
rect 20605 92807 20639 92835
rect 20667 92807 20701 92835
rect 20729 92807 20763 92835
rect 20791 92807 20839 92835
rect 20529 92773 20839 92807
rect 20529 92745 20577 92773
rect 20605 92745 20639 92773
rect 20667 92745 20701 92773
rect 20729 92745 20763 92773
rect 20791 92745 20839 92773
rect 13389 86931 13437 86959
rect 13465 86931 13499 86959
rect 13527 86931 13561 86959
rect 13589 86931 13623 86959
rect 13651 86931 13699 86959
rect 13389 86897 13699 86931
rect 13389 86869 13437 86897
rect 13465 86869 13499 86897
rect 13527 86869 13561 86897
rect 13589 86869 13623 86897
rect 13651 86869 13699 86897
rect 13389 86835 13699 86869
rect 13389 86807 13437 86835
rect 13465 86807 13499 86835
rect 13527 86807 13561 86835
rect 13589 86807 13623 86835
rect 13651 86807 13699 86835
rect 13389 86773 13699 86807
rect 13389 86745 13437 86773
rect 13465 86745 13499 86773
rect 13527 86745 13561 86773
rect 13589 86745 13623 86773
rect 13651 86745 13699 86773
rect 13389 77959 13699 86745
rect 17224 83959 17384 83976
rect 17224 83931 17259 83959
rect 17287 83931 17321 83959
rect 17349 83931 17384 83959
rect 17224 83897 17384 83931
rect 17224 83869 17259 83897
rect 17287 83869 17321 83897
rect 17349 83869 17384 83897
rect 17224 83835 17384 83869
rect 17224 83807 17259 83835
rect 17287 83807 17321 83835
rect 17349 83807 17384 83835
rect 17224 83773 17384 83807
rect 17224 83745 17259 83773
rect 17287 83745 17321 83773
rect 17349 83745 17384 83773
rect 17224 83728 17384 83745
rect 20529 83959 20839 92745
rect 20529 83931 20577 83959
rect 20605 83931 20639 83959
rect 20667 83931 20701 83959
rect 20729 83931 20763 83959
rect 20791 83931 20839 83959
rect 20529 83897 20839 83931
rect 20529 83869 20577 83897
rect 20605 83869 20639 83897
rect 20667 83869 20701 83897
rect 20729 83869 20763 83897
rect 20791 83869 20839 83897
rect 20529 83835 20839 83869
rect 20529 83807 20577 83835
rect 20605 83807 20639 83835
rect 20667 83807 20701 83835
rect 20729 83807 20763 83835
rect 20791 83807 20839 83835
rect 20529 83773 20839 83807
rect 20529 83745 20577 83773
rect 20605 83745 20639 83773
rect 20667 83745 20701 83773
rect 20729 83745 20763 83773
rect 20791 83745 20839 83773
rect 13389 77931 13437 77959
rect 13465 77931 13499 77959
rect 13527 77931 13561 77959
rect 13589 77931 13623 77959
rect 13651 77931 13699 77959
rect 13389 77897 13699 77931
rect 13389 77869 13437 77897
rect 13465 77869 13499 77897
rect 13527 77869 13561 77897
rect 13589 77869 13623 77897
rect 13651 77869 13699 77897
rect 13389 77835 13699 77869
rect 13389 77807 13437 77835
rect 13465 77807 13499 77835
rect 13527 77807 13561 77835
rect 13589 77807 13623 77835
rect 13651 77807 13699 77835
rect 13389 77773 13699 77807
rect 13389 77745 13437 77773
rect 13465 77745 13499 77773
rect 13527 77745 13561 77773
rect 13589 77745 13623 77773
rect 13651 77745 13699 77773
rect 13389 68959 13699 77745
rect 17224 74959 17384 74976
rect 17224 74931 17259 74959
rect 17287 74931 17321 74959
rect 17349 74931 17384 74959
rect 17224 74897 17384 74931
rect 17224 74869 17259 74897
rect 17287 74869 17321 74897
rect 17349 74869 17384 74897
rect 17224 74835 17384 74869
rect 17224 74807 17259 74835
rect 17287 74807 17321 74835
rect 17349 74807 17384 74835
rect 17224 74773 17384 74807
rect 17224 74745 17259 74773
rect 17287 74745 17321 74773
rect 17349 74745 17384 74773
rect 17224 74728 17384 74745
rect 20529 74959 20839 83745
rect 20529 74931 20577 74959
rect 20605 74931 20639 74959
rect 20667 74931 20701 74959
rect 20729 74931 20763 74959
rect 20791 74931 20839 74959
rect 20529 74897 20839 74931
rect 20529 74869 20577 74897
rect 20605 74869 20639 74897
rect 20667 74869 20701 74897
rect 20729 74869 20763 74897
rect 20791 74869 20839 74897
rect 20529 74835 20839 74869
rect 20529 74807 20577 74835
rect 20605 74807 20639 74835
rect 20667 74807 20701 74835
rect 20729 74807 20763 74835
rect 20791 74807 20839 74835
rect 20529 74773 20839 74807
rect 20529 74745 20577 74773
rect 20605 74745 20639 74773
rect 20667 74745 20701 74773
rect 20729 74745 20763 74773
rect 20791 74745 20839 74773
rect 13389 68931 13437 68959
rect 13465 68931 13499 68959
rect 13527 68931 13561 68959
rect 13589 68931 13623 68959
rect 13651 68931 13699 68959
rect 13389 68897 13699 68931
rect 13389 68869 13437 68897
rect 13465 68869 13499 68897
rect 13527 68869 13561 68897
rect 13589 68869 13623 68897
rect 13651 68869 13699 68897
rect 13389 68835 13699 68869
rect 13389 68807 13437 68835
rect 13465 68807 13499 68835
rect 13527 68807 13561 68835
rect 13589 68807 13623 68835
rect 13651 68807 13699 68835
rect 13389 68773 13699 68807
rect 13389 68745 13437 68773
rect 13465 68745 13499 68773
rect 13527 68745 13561 68773
rect 13589 68745 13623 68773
rect 13651 68745 13699 68773
rect 13389 59959 13699 68745
rect 17224 65959 17384 65976
rect 17224 65931 17259 65959
rect 17287 65931 17321 65959
rect 17349 65931 17384 65959
rect 17224 65897 17384 65931
rect 17224 65869 17259 65897
rect 17287 65869 17321 65897
rect 17349 65869 17384 65897
rect 17224 65835 17384 65869
rect 17224 65807 17259 65835
rect 17287 65807 17321 65835
rect 17349 65807 17384 65835
rect 17224 65773 17384 65807
rect 17224 65745 17259 65773
rect 17287 65745 17321 65773
rect 17349 65745 17384 65773
rect 17224 65728 17384 65745
rect 20529 65959 20839 74745
rect 20529 65931 20577 65959
rect 20605 65931 20639 65959
rect 20667 65931 20701 65959
rect 20729 65931 20763 65959
rect 20791 65931 20839 65959
rect 20529 65897 20839 65931
rect 20529 65869 20577 65897
rect 20605 65869 20639 65897
rect 20667 65869 20701 65897
rect 20729 65869 20763 65897
rect 20791 65869 20839 65897
rect 20529 65835 20839 65869
rect 20529 65807 20577 65835
rect 20605 65807 20639 65835
rect 20667 65807 20701 65835
rect 20729 65807 20763 65835
rect 20791 65807 20839 65835
rect 20529 65773 20839 65807
rect 20529 65745 20577 65773
rect 20605 65745 20639 65773
rect 20667 65745 20701 65773
rect 20729 65745 20763 65773
rect 20791 65745 20839 65773
rect 13389 59931 13437 59959
rect 13465 59931 13499 59959
rect 13527 59931 13561 59959
rect 13589 59931 13623 59959
rect 13651 59931 13699 59959
rect 13389 59897 13699 59931
rect 13389 59869 13437 59897
rect 13465 59869 13499 59897
rect 13527 59869 13561 59897
rect 13589 59869 13623 59897
rect 13651 59869 13699 59897
rect 13389 59835 13699 59869
rect 13389 59807 13437 59835
rect 13465 59807 13499 59835
rect 13527 59807 13561 59835
rect 13589 59807 13623 59835
rect 13651 59807 13699 59835
rect 13389 59773 13699 59807
rect 13389 59745 13437 59773
rect 13465 59745 13499 59773
rect 13527 59745 13561 59773
rect 13589 59745 13623 59773
rect 13651 59745 13699 59773
rect 13389 50959 13699 59745
rect 17224 56959 17384 56976
rect 17224 56931 17259 56959
rect 17287 56931 17321 56959
rect 17349 56931 17384 56959
rect 17224 56897 17384 56931
rect 17224 56869 17259 56897
rect 17287 56869 17321 56897
rect 17349 56869 17384 56897
rect 17224 56835 17384 56869
rect 17224 56807 17259 56835
rect 17287 56807 17321 56835
rect 17349 56807 17384 56835
rect 17224 56773 17384 56807
rect 17224 56745 17259 56773
rect 17287 56745 17321 56773
rect 17349 56745 17384 56773
rect 17224 56728 17384 56745
rect 20529 56959 20839 65745
rect 20529 56931 20577 56959
rect 20605 56931 20639 56959
rect 20667 56931 20701 56959
rect 20729 56931 20763 56959
rect 20791 56931 20839 56959
rect 20529 56897 20839 56931
rect 20529 56869 20577 56897
rect 20605 56869 20639 56897
rect 20667 56869 20701 56897
rect 20729 56869 20763 56897
rect 20791 56869 20839 56897
rect 20529 56835 20839 56869
rect 20529 56807 20577 56835
rect 20605 56807 20639 56835
rect 20667 56807 20701 56835
rect 20729 56807 20763 56835
rect 20791 56807 20839 56835
rect 20529 56773 20839 56807
rect 20529 56745 20577 56773
rect 20605 56745 20639 56773
rect 20667 56745 20701 56773
rect 20729 56745 20763 56773
rect 20791 56745 20839 56773
rect 13389 50931 13437 50959
rect 13465 50931 13499 50959
rect 13527 50931 13561 50959
rect 13589 50931 13623 50959
rect 13651 50931 13699 50959
rect 13389 50897 13699 50931
rect 13389 50869 13437 50897
rect 13465 50869 13499 50897
rect 13527 50869 13561 50897
rect 13589 50869 13623 50897
rect 13651 50869 13699 50897
rect 13389 50835 13699 50869
rect 13389 50807 13437 50835
rect 13465 50807 13499 50835
rect 13527 50807 13561 50835
rect 13589 50807 13623 50835
rect 13651 50807 13699 50835
rect 13389 50773 13699 50807
rect 13389 50745 13437 50773
rect 13465 50745 13499 50773
rect 13527 50745 13561 50773
rect 13589 50745 13623 50773
rect 13651 50745 13699 50773
rect 13389 41959 13699 50745
rect 17224 47959 17384 47976
rect 17224 47931 17259 47959
rect 17287 47931 17321 47959
rect 17349 47931 17384 47959
rect 17224 47897 17384 47931
rect 17224 47869 17259 47897
rect 17287 47869 17321 47897
rect 17349 47869 17384 47897
rect 17224 47835 17384 47869
rect 17224 47807 17259 47835
rect 17287 47807 17321 47835
rect 17349 47807 17384 47835
rect 17224 47773 17384 47807
rect 17224 47745 17259 47773
rect 17287 47745 17321 47773
rect 17349 47745 17384 47773
rect 17224 47728 17384 47745
rect 20529 47959 20839 56745
rect 20529 47931 20577 47959
rect 20605 47931 20639 47959
rect 20667 47931 20701 47959
rect 20729 47931 20763 47959
rect 20791 47931 20839 47959
rect 20529 47897 20839 47931
rect 20529 47869 20577 47897
rect 20605 47869 20639 47897
rect 20667 47869 20701 47897
rect 20729 47869 20763 47897
rect 20791 47869 20839 47897
rect 20529 47835 20839 47869
rect 20529 47807 20577 47835
rect 20605 47807 20639 47835
rect 20667 47807 20701 47835
rect 20729 47807 20763 47835
rect 20791 47807 20839 47835
rect 20529 47773 20839 47807
rect 20529 47745 20577 47773
rect 20605 47745 20639 47773
rect 20667 47745 20701 47773
rect 20729 47745 20763 47773
rect 20791 47745 20839 47773
rect 13389 41931 13437 41959
rect 13465 41931 13499 41959
rect 13527 41931 13561 41959
rect 13589 41931 13623 41959
rect 13651 41931 13699 41959
rect 13389 41897 13699 41931
rect 13389 41869 13437 41897
rect 13465 41869 13499 41897
rect 13527 41869 13561 41897
rect 13589 41869 13623 41897
rect 13651 41869 13699 41897
rect 13389 41835 13699 41869
rect 13389 41807 13437 41835
rect 13465 41807 13499 41835
rect 13527 41807 13561 41835
rect 13589 41807 13623 41835
rect 13651 41807 13699 41835
rect 13389 41773 13699 41807
rect 13389 41745 13437 41773
rect 13465 41745 13499 41773
rect 13527 41745 13561 41773
rect 13589 41745 13623 41773
rect 13651 41745 13699 41773
rect 13389 32959 13699 41745
rect 17224 38959 17384 38976
rect 17224 38931 17259 38959
rect 17287 38931 17321 38959
rect 17349 38931 17384 38959
rect 17224 38897 17384 38931
rect 17224 38869 17259 38897
rect 17287 38869 17321 38897
rect 17349 38869 17384 38897
rect 17224 38835 17384 38869
rect 17224 38807 17259 38835
rect 17287 38807 17321 38835
rect 17349 38807 17384 38835
rect 17224 38773 17384 38807
rect 17224 38745 17259 38773
rect 17287 38745 17321 38773
rect 17349 38745 17384 38773
rect 17224 38728 17384 38745
rect 20529 38959 20839 47745
rect 20529 38931 20577 38959
rect 20605 38931 20639 38959
rect 20667 38931 20701 38959
rect 20729 38931 20763 38959
rect 20791 38931 20839 38959
rect 20529 38897 20839 38931
rect 20529 38869 20577 38897
rect 20605 38869 20639 38897
rect 20667 38869 20701 38897
rect 20729 38869 20763 38897
rect 20791 38869 20839 38897
rect 20529 38835 20839 38869
rect 20529 38807 20577 38835
rect 20605 38807 20639 38835
rect 20667 38807 20701 38835
rect 20729 38807 20763 38835
rect 20791 38807 20839 38835
rect 20529 38773 20839 38807
rect 20529 38745 20577 38773
rect 20605 38745 20639 38773
rect 20667 38745 20701 38773
rect 20729 38745 20763 38773
rect 20791 38745 20839 38773
rect 13389 32931 13437 32959
rect 13465 32931 13499 32959
rect 13527 32931 13561 32959
rect 13589 32931 13623 32959
rect 13651 32931 13699 32959
rect 13389 32897 13699 32931
rect 13389 32869 13437 32897
rect 13465 32869 13499 32897
rect 13527 32869 13561 32897
rect 13589 32869 13623 32897
rect 13651 32869 13699 32897
rect 13389 32835 13699 32869
rect 13389 32807 13437 32835
rect 13465 32807 13499 32835
rect 13527 32807 13561 32835
rect 13589 32807 13623 32835
rect 13651 32807 13699 32835
rect 13389 32773 13699 32807
rect 13389 32745 13437 32773
rect 13465 32745 13499 32773
rect 13527 32745 13561 32773
rect 13589 32745 13623 32773
rect 13651 32745 13699 32773
rect 13389 23959 13699 32745
rect 17224 29959 17384 29976
rect 17224 29931 17259 29959
rect 17287 29931 17321 29959
rect 17349 29931 17384 29959
rect 17224 29897 17384 29931
rect 17224 29869 17259 29897
rect 17287 29869 17321 29897
rect 17349 29869 17384 29897
rect 17224 29835 17384 29869
rect 17224 29807 17259 29835
rect 17287 29807 17321 29835
rect 17349 29807 17384 29835
rect 17224 29773 17384 29807
rect 17224 29745 17259 29773
rect 17287 29745 17321 29773
rect 17349 29745 17384 29773
rect 17224 29728 17384 29745
rect 20529 29959 20839 38745
rect 20529 29931 20577 29959
rect 20605 29931 20639 29959
rect 20667 29931 20701 29959
rect 20729 29931 20763 29959
rect 20791 29931 20839 29959
rect 20529 29897 20839 29931
rect 20529 29869 20577 29897
rect 20605 29869 20639 29897
rect 20667 29869 20701 29897
rect 20729 29869 20763 29897
rect 20791 29869 20839 29897
rect 20529 29835 20839 29869
rect 20529 29807 20577 29835
rect 20605 29807 20639 29835
rect 20667 29807 20701 29835
rect 20729 29807 20763 29835
rect 20791 29807 20839 29835
rect 20529 29773 20839 29807
rect 20529 29745 20577 29773
rect 20605 29745 20639 29773
rect 20667 29745 20701 29773
rect 20729 29745 20763 29773
rect 20791 29745 20839 29773
rect 13389 23931 13437 23959
rect 13465 23931 13499 23959
rect 13527 23931 13561 23959
rect 13589 23931 13623 23959
rect 13651 23931 13699 23959
rect 13389 23897 13699 23931
rect 13389 23869 13437 23897
rect 13465 23869 13499 23897
rect 13527 23869 13561 23897
rect 13589 23869 13623 23897
rect 13651 23869 13699 23897
rect 13389 23835 13699 23869
rect 13389 23807 13437 23835
rect 13465 23807 13499 23835
rect 13527 23807 13561 23835
rect 13589 23807 13623 23835
rect 13651 23807 13699 23835
rect 13389 23773 13699 23807
rect 13389 23745 13437 23773
rect 13465 23745 13499 23773
rect 13527 23745 13561 23773
rect 13589 23745 13623 23773
rect 13651 23745 13699 23773
rect 13389 14959 13699 23745
rect 17224 20959 17384 20976
rect 17224 20931 17259 20959
rect 17287 20931 17321 20959
rect 17349 20931 17384 20959
rect 17224 20897 17384 20931
rect 17224 20869 17259 20897
rect 17287 20869 17321 20897
rect 17349 20869 17384 20897
rect 17224 20835 17384 20869
rect 17224 20807 17259 20835
rect 17287 20807 17321 20835
rect 17349 20807 17384 20835
rect 17224 20773 17384 20807
rect 17224 20745 17259 20773
rect 17287 20745 17321 20773
rect 17349 20745 17384 20773
rect 17224 20728 17384 20745
rect 20529 20959 20839 29745
rect 20529 20931 20577 20959
rect 20605 20931 20639 20959
rect 20667 20931 20701 20959
rect 20729 20931 20763 20959
rect 20791 20931 20839 20959
rect 20529 20897 20839 20931
rect 20529 20869 20577 20897
rect 20605 20869 20639 20897
rect 20667 20869 20701 20897
rect 20729 20869 20763 20897
rect 20791 20869 20839 20897
rect 20529 20835 20839 20869
rect 20529 20807 20577 20835
rect 20605 20807 20639 20835
rect 20667 20807 20701 20835
rect 20729 20807 20763 20835
rect 20791 20807 20839 20835
rect 20529 20773 20839 20807
rect 20529 20745 20577 20773
rect 20605 20745 20639 20773
rect 20667 20745 20701 20773
rect 20729 20745 20763 20773
rect 20791 20745 20839 20773
rect 13389 14931 13437 14959
rect 13465 14931 13499 14959
rect 13527 14931 13561 14959
rect 13589 14931 13623 14959
rect 13651 14931 13699 14959
rect 13389 14897 13699 14931
rect 13389 14869 13437 14897
rect 13465 14869 13499 14897
rect 13527 14869 13561 14897
rect 13589 14869 13623 14897
rect 13651 14869 13699 14897
rect 13389 14835 13699 14869
rect 13389 14807 13437 14835
rect 13465 14807 13499 14835
rect 13527 14807 13561 14835
rect 13589 14807 13623 14835
rect 13651 14807 13699 14835
rect 13389 14773 13699 14807
rect 13389 14745 13437 14773
rect 13465 14745 13499 14773
rect 13527 14745 13561 14773
rect 13589 14745 13623 14773
rect 13651 14745 13699 14773
rect 13389 5959 13699 14745
rect 13389 5931 13437 5959
rect 13465 5931 13499 5959
rect 13527 5931 13561 5959
rect 13589 5931 13623 5959
rect 13651 5931 13699 5959
rect 13389 5897 13699 5931
rect 13389 5869 13437 5897
rect 13465 5869 13499 5897
rect 13527 5869 13561 5897
rect 13589 5869 13623 5897
rect 13651 5869 13699 5897
rect 13389 5835 13699 5869
rect 13389 5807 13437 5835
rect 13465 5807 13499 5835
rect 13527 5807 13561 5835
rect 13589 5807 13623 5835
rect 13651 5807 13699 5835
rect 13389 5773 13699 5807
rect 13389 5745 13437 5773
rect 13465 5745 13499 5773
rect 13527 5745 13561 5773
rect 13589 5745 13623 5773
rect 13651 5745 13699 5773
rect 13389 424 13699 5745
rect 13389 396 13437 424
rect 13465 396 13499 424
rect 13527 396 13561 424
rect 13589 396 13623 424
rect 13651 396 13699 424
rect 13389 362 13699 396
rect 13389 334 13437 362
rect 13465 334 13499 362
rect 13527 334 13561 362
rect 13589 334 13623 362
rect 13651 334 13699 362
rect 13389 300 13699 334
rect 13389 272 13437 300
rect 13465 272 13499 300
rect 13527 272 13561 300
rect 13589 272 13623 300
rect 13651 272 13699 300
rect 13389 238 13699 272
rect 13389 210 13437 238
rect 13465 210 13499 238
rect 13527 210 13561 238
rect 13589 210 13623 238
rect 13651 210 13699 238
rect 13389 162 13699 210
rect 20529 11959 20839 20745
rect 20529 11931 20577 11959
rect 20605 11931 20639 11959
rect 20667 11931 20701 11959
rect 20729 11931 20763 11959
rect 20791 11931 20839 11959
rect 20529 11897 20839 11931
rect 20529 11869 20577 11897
rect 20605 11869 20639 11897
rect 20667 11869 20701 11897
rect 20729 11869 20763 11897
rect 20791 11869 20839 11897
rect 20529 11835 20839 11869
rect 20529 11807 20577 11835
rect 20605 11807 20639 11835
rect 20667 11807 20701 11835
rect 20729 11807 20763 11835
rect 20791 11807 20839 11835
rect 20529 11773 20839 11807
rect 20529 11745 20577 11773
rect 20605 11745 20639 11773
rect 20667 11745 20701 11773
rect 20729 11745 20763 11773
rect 20791 11745 20839 11773
rect 20529 2959 20839 11745
rect 20529 2931 20577 2959
rect 20605 2931 20639 2959
rect 20667 2931 20701 2959
rect 20729 2931 20763 2959
rect 20791 2931 20839 2959
rect 20529 2897 20839 2931
rect 20529 2869 20577 2897
rect 20605 2869 20639 2897
rect 20667 2869 20701 2897
rect 20729 2869 20763 2897
rect 20791 2869 20839 2897
rect 20529 2835 20839 2869
rect 20529 2807 20577 2835
rect 20605 2807 20639 2835
rect 20667 2807 20701 2835
rect 20729 2807 20763 2835
rect 20791 2807 20839 2835
rect 20529 2773 20839 2807
rect 20529 2745 20577 2773
rect 20605 2745 20639 2773
rect 20667 2745 20701 2773
rect 20729 2745 20763 2773
rect 20791 2745 20839 2773
rect 20529 904 20839 2745
rect 20529 876 20577 904
rect 20605 876 20639 904
rect 20667 876 20701 904
rect 20729 876 20763 904
rect 20791 876 20839 904
rect 20529 842 20839 876
rect 20529 814 20577 842
rect 20605 814 20639 842
rect 20667 814 20701 842
rect 20729 814 20763 842
rect 20791 814 20839 842
rect 20529 780 20839 814
rect 20529 752 20577 780
rect 20605 752 20639 780
rect 20667 752 20701 780
rect 20729 752 20763 780
rect 20791 752 20839 780
rect 20529 718 20839 752
rect 20529 690 20577 718
rect 20605 690 20639 718
rect 20667 690 20701 718
rect 20729 690 20763 718
rect 20791 690 20839 718
rect 20529 162 20839 690
rect 22389 299670 22699 299718
rect 22389 299642 22437 299670
rect 22465 299642 22499 299670
rect 22527 299642 22561 299670
rect 22589 299642 22623 299670
rect 22651 299642 22699 299670
rect 22389 299608 22699 299642
rect 22389 299580 22437 299608
rect 22465 299580 22499 299608
rect 22527 299580 22561 299608
rect 22589 299580 22623 299608
rect 22651 299580 22699 299608
rect 22389 299546 22699 299580
rect 22389 299518 22437 299546
rect 22465 299518 22499 299546
rect 22527 299518 22561 299546
rect 22589 299518 22623 299546
rect 22651 299518 22699 299546
rect 22389 299484 22699 299518
rect 22389 299456 22437 299484
rect 22465 299456 22499 299484
rect 22527 299456 22561 299484
rect 22589 299456 22623 299484
rect 22651 299456 22699 299484
rect 22389 293959 22699 299456
rect 22389 293931 22437 293959
rect 22465 293931 22499 293959
rect 22527 293931 22561 293959
rect 22589 293931 22623 293959
rect 22651 293931 22699 293959
rect 22389 293897 22699 293931
rect 22389 293869 22437 293897
rect 22465 293869 22499 293897
rect 22527 293869 22561 293897
rect 22589 293869 22623 293897
rect 22651 293869 22699 293897
rect 22389 293835 22699 293869
rect 22389 293807 22437 293835
rect 22465 293807 22499 293835
rect 22527 293807 22561 293835
rect 22589 293807 22623 293835
rect 22651 293807 22699 293835
rect 22389 293773 22699 293807
rect 22389 293745 22437 293773
rect 22465 293745 22499 293773
rect 22527 293745 22561 293773
rect 22589 293745 22623 293773
rect 22651 293745 22699 293773
rect 22389 284959 22699 293745
rect 22389 284931 22437 284959
rect 22465 284931 22499 284959
rect 22527 284931 22561 284959
rect 22589 284931 22623 284959
rect 22651 284931 22699 284959
rect 22389 284897 22699 284931
rect 22389 284869 22437 284897
rect 22465 284869 22499 284897
rect 22527 284869 22561 284897
rect 22589 284869 22623 284897
rect 22651 284869 22699 284897
rect 22389 284835 22699 284869
rect 22389 284807 22437 284835
rect 22465 284807 22499 284835
rect 22527 284807 22561 284835
rect 22589 284807 22623 284835
rect 22651 284807 22699 284835
rect 22389 284773 22699 284807
rect 22389 284745 22437 284773
rect 22465 284745 22499 284773
rect 22527 284745 22561 284773
rect 22589 284745 22623 284773
rect 22651 284745 22699 284773
rect 22389 275959 22699 284745
rect 22389 275931 22437 275959
rect 22465 275931 22499 275959
rect 22527 275931 22561 275959
rect 22589 275931 22623 275959
rect 22651 275931 22699 275959
rect 22389 275897 22699 275931
rect 22389 275869 22437 275897
rect 22465 275869 22499 275897
rect 22527 275869 22561 275897
rect 22589 275869 22623 275897
rect 22651 275869 22699 275897
rect 22389 275835 22699 275869
rect 22389 275807 22437 275835
rect 22465 275807 22499 275835
rect 22527 275807 22561 275835
rect 22589 275807 22623 275835
rect 22651 275807 22699 275835
rect 22389 275773 22699 275807
rect 22389 275745 22437 275773
rect 22465 275745 22499 275773
rect 22527 275745 22561 275773
rect 22589 275745 22623 275773
rect 22651 275745 22699 275773
rect 22389 266959 22699 275745
rect 22389 266931 22437 266959
rect 22465 266931 22499 266959
rect 22527 266931 22561 266959
rect 22589 266931 22623 266959
rect 22651 266931 22699 266959
rect 22389 266897 22699 266931
rect 22389 266869 22437 266897
rect 22465 266869 22499 266897
rect 22527 266869 22561 266897
rect 22589 266869 22623 266897
rect 22651 266869 22699 266897
rect 22389 266835 22699 266869
rect 22389 266807 22437 266835
rect 22465 266807 22499 266835
rect 22527 266807 22561 266835
rect 22589 266807 22623 266835
rect 22651 266807 22699 266835
rect 22389 266773 22699 266807
rect 22389 266745 22437 266773
rect 22465 266745 22499 266773
rect 22527 266745 22561 266773
rect 22589 266745 22623 266773
rect 22651 266745 22699 266773
rect 22389 257959 22699 266745
rect 22389 257931 22437 257959
rect 22465 257931 22499 257959
rect 22527 257931 22561 257959
rect 22589 257931 22623 257959
rect 22651 257931 22699 257959
rect 22389 257897 22699 257931
rect 22389 257869 22437 257897
rect 22465 257869 22499 257897
rect 22527 257869 22561 257897
rect 22589 257869 22623 257897
rect 22651 257869 22699 257897
rect 22389 257835 22699 257869
rect 22389 257807 22437 257835
rect 22465 257807 22499 257835
rect 22527 257807 22561 257835
rect 22589 257807 22623 257835
rect 22651 257807 22699 257835
rect 22389 257773 22699 257807
rect 22389 257745 22437 257773
rect 22465 257745 22499 257773
rect 22527 257745 22561 257773
rect 22589 257745 22623 257773
rect 22651 257745 22699 257773
rect 22389 248959 22699 257745
rect 29529 299190 29839 299718
rect 29529 299162 29577 299190
rect 29605 299162 29639 299190
rect 29667 299162 29701 299190
rect 29729 299162 29763 299190
rect 29791 299162 29839 299190
rect 29529 299128 29839 299162
rect 29529 299100 29577 299128
rect 29605 299100 29639 299128
rect 29667 299100 29701 299128
rect 29729 299100 29763 299128
rect 29791 299100 29839 299128
rect 29529 299066 29839 299100
rect 29529 299038 29577 299066
rect 29605 299038 29639 299066
rect 29667 299038 29701 299066
rect 29729 299038 29763 299066
rect 29791 299038 29839 299066
rect 29529 299004 29839 299038
rect 29529 298976 29577 299004
rect 29605 298976 29639 299004
rect 29667 298976 29701 299004
rect 29729 298976 29763 299004
rect 29791 298976 29839 299004
rect 29529 290959 29839 298976
rect 29529 290931 29577 290959
rect 29605 290931 29639 290959
rect 29667 290931 29701 290959
rect 29729 290931 29763 290959
rect 29791 290931 29839 290959
rect 29529 290897 29839 290931
rect 29529 290869 29577 290897
rect 29605 290869 29639 290897
rect 29667 290869 29701 290897
rect 29729 290869 29763 290897
rect 29791 290869 29839 290897
rect 29529 290835 29839 290869
rect 29529 290807 29577 290835
rect 29605 290807 29639 290835
rect 29667 290807 29701 290835
rect 29729 290807 29763 290835
rect 29791 290807 29839 290835
rect 29529 290773 29839 290807
rect 29529 290745 29577 290773
rect 29605 290745 29639 290773
rect 29667 290745 29701 290773
rect 29729 290745 29763 290773
rect 29791 290745 29839 290773
rect 29529 281959 29839 290745
rect 29529 281931 29577 281959
rect 29605 281931 29639 281959
rect 29667 281931 29701 281959
rect 29729 281931 29763 281959
rect 29791 281931 29839 281959
rect 29529 281897 29839 281931
rect 29529 281869 29577 281897
rect 29605 281869 29639 281897
rect 29667 281869 29701 281897
rect 29729 281869 29763 281897
rect 29791 281869 29839 281897
rect 29529 281835 29839 281869
rect 29529 281807 29577 281835
rect 29605 281807 29639 281835
rect 29667 281807 29701 281835
rect 29729 281807 29763 281835
rect 29791 281807 29839 281835
rect 29529 281773 29839 281807
rect 29529 281745 29577 281773
rect 29605 281745 29639 281773
rect 29667 281745 29701 281773
rect 29729 281745 29763 281773
rect 29791 281745 29839 281773
rect 29529 272959 29839 281745
rect 29529 272931 29577 272959
rect 29605 272931 29639 272959
rect 29667 272931 29701 272959
rect 29729 272931 29763 272959
rect 29791 272931 29839 272959
rect 29529 272897 29839 272931
rect 29529 272869 29577 272897
rect 29605 272869 29639 272897
rect 29667 272869 29701 272897
rect 29729 272869 29763 272897
rect 29791 272869 29839 272897
rect 29529 272835 29839 272869
rect 29529 272807 29577 272835
rect 29605 272807 29639 272835
rect 29667 272807 29701 272835
rect 29729 272807 29763 272835
rect 29791 272807 29839 272835
rect 29529 272773 29839 272807
rect 29529 272745 29577 272773
rect 29605 272745 29639 272773
rect 29667 272745 29701 272773
rect 29729 272745 29763 272773
rect 29791 272745 29839 272773
rect 29529 263959 29839 272745
rect 29529 263931 29577 263959
rect 29605 263931 29639 263959
rect 29667 263931 29701 263959
rect 29729 263931 29763 263959
rect 29791 263931 29839 263959
rect 29529 263897 29839 263931
rect 29529 263869 29577 263897
rect 29605 263869 29639 263897
rect 29667 263869 29701 263897
rect 29729 263869 29763 263897
rect 29791 263869 29839 263897
rect 29529 263835 29839 263869
rect 29529 263807 29577 263835
rect 29605 263807 29639 263835
rect 29667 263807 29701 263835
rect 29729 263807 29763 263835
rect 29791 263807 29839 263835
rect 29529 263773 29839 263807
rect 29529 263745 29577 263773
rect 29605 263745 29639 263773
rect 29667 263745 29701 263773
rect 29729 263745 29763 263773
rect 29791 263745 29839 263773
rect 29529 254959 29839 263745
rect 29529 254931 29577 254959
rect 29605 254931 29639 254959
rect 29667 254931 29701 254959
rect 29729 254931 29763 254959
rect 29791 254931 29839 254959
rect 29529 254897 29839 254931
rect 29529 254869 29577 254897
rect 29605 254869 29639 254897
rect 29667 254869 29701 254897
rect 29729 254869 29763 254897
rect 29791 254869 29839 254897
rect 29529 254835 29839 254869
rect 29529 254807 29577 254835
rect 29605 254807 29639 254835
rect 29667 254807 29701 254835
rect 29729 254807 29763 254835
rect 29791 254807 29839 254835
rect 29529 254773 29839 254807
rect 29529 254745 29577 254773
rect 29605 254745 29639 254773
rect 29667 254745 29701 254773
rect 29729 254745 29763 254773
rect 29791 254745 29839 254773
rect 22389 248931 22437 248959
rect 22465 248931 22499 248959
rect 22527 248931 22561 248959
rect 22589 248931 22623 248959
rect 22651 248931 22699 248959
rect 22389 248897 22699 248931
rect 22389 248869 22437 248897
rect 22465 248869 22499 248897
rect 22527 248869 22561 248897
rect 22589 248869 22623 248897
rect 22651 248869 22699 248897
rect 22389 248835 22699 248869
rect 22389 248807 22437 248835
rect 22465 248807 22499 248835
rect 22527 248807 22561 248835
rect 22589 248807 22623 248835
rect 22651 248807 22699 248835
rect 22389 248773 22699 248807
rect 22389 248745 22437 248773
rect 22465 248745 22499 248773
rect 22527 248745 22561 248773
rect 22589 248745 22623 248773
rect 22651 248745 22699 248773
rect 22389 239959 22699 248745
rect 24904 248959 25064 248976
rect 24904 248931 24939 248959
rect 24967 248931 25001 248959
rect 25029 248931 25064 248959
rect 24904 248897 25064 248931
rect 24904 248869 24939 248897
rect 24967 248869 25001 248897
rect 25029 248869 25064 248897
rect 24904 248835 25064 248869
rect 24904 248807 24939 248835
rect 24967 248807 25001 248835
rect 25029 248807 25064 248835
rect 24904 248773 25064 248807
rect 24904 248745 24939 248773
rect 24967 248745 25001 248773
rect 25029 248745 25064 248773
rect 24904 248728 25064 248745
rect 29529 245959 29839 254745
rect 29529 245931 29577 245959
rect 29605 245931 29639 245959
rect 29667 245931 29701 245959
rect 29729 245931 29763 245959
rect 29791 245931 29839 245959
rect 29529 245897 29839 245931
rect 29529 245869 29577 245897
rect 29605 245869 29639 245897
rect 29667 245869 29701 245897
rect 29729 245869 29763 245897
rect 29791 245869 29839 245897
rect 29529 245835 29839 245869
rect 29529 245807 29577 245835
rect 29605 245807 29639 245835
rect 29667 245807 29701 245835
rect 29729 245807 29763 245835
rect 29791 245807 29839 245835
rect 29529 245773 29839 245807
rect 29529 245745 29577 245773
rect 29605 245745 29639 245773
rect 29667 245745 29701 245773
rect 29729 245745 29763 245773
rect 29791 245745 29839 245773
rect 22389 239931 22437 239959
rect 22465 239931 22499 239959
rect 22527 239931 22561 239959
rect 22589 239931 22623 239959
rect 22651 239931 22699 239959
rect 22389 239897 22699 239931
rect 22389 239869 22437 239897
rect 22465 239869 22499 239897
rect 22527 239869 22561 239897
rect 22589 239869 22623 239897
rect 22651 239869 22699 239897
rect 22389 239835 22699 239869
rect 22389 239807 22437 239835
rect 22465 239807 22499 239835
rect 22527 239807 22561 239835
rect 22589 239807 22623 239835
rect 22651 239807 22699 239835
rect 22389 239773 22699 239807
rect 22389 239745 22437 239773
rect 22465 239745 22499 239773
rect 22527 239745 22561 239773
rect 22589 239745 22623 239773
rect 22651 239745 22699 239773
rect 22389 230959 22699 239745
rect 24904 239959 25064 239976
rect 24904 239931 24939 239959
rect 24967 239931 25001 239959
rect 25029 239931 25064 239959
rect 24904 239897 25064 239931
rect 24904 239869 24939 239897
rect 24967 239869 25001 239897
rect 25029 239869 25064 239897
rect 24904 239835 25064 239869
rect 24904 239807 24939 239835
rect 24967 239807 25001 239835
rect 25029 239807 25064 239835
rect 24904 239773 25064 239807
rect 24904 239745 24939 239773
rect 24967 239745 25001 239773
rect 25029 239745 25064 239773
rect 24904 239728 25064 239745
rect 29529 236959 29839 245745
rect 29529 236931 29577 236959
rect 29605 236931 29639 236959
rect 29667 236931 29701 236959
rect 29729 236931 29763 236959
rect 29791 236931 29839 236959
rect 29529 236897 29839 236931
rect 29529 236869 29577 236897
rect 29605 236869 29639 236897
rect 29667 236869 29701 236897
rect 29729 236869 29763 236897
rect 29791 236869 29839 236897
rect 29529 236835 29839 236869
rect 29529 236807 29577 236835
rect 29605 236807 29639 236835
rect 29667 236807 29701 236835
rect 29729 236807 29763 236835
rect 29791 236807 29839 236835
rect 29529 236773 29839 236807
rect 29529 236745 29577 236773
rect 29605 236745 29639 236773
rect 29667 236745 29701 236773
rect 29729 236745 29763 236773
rect 29791 236745 29839 236773
rect 22389 230931 22437 230959
rect 22465 230931 22499 230959
rect 22527 230931 22561 230959
rect 22589 230931 22623 230959
rect 22651 230931 22699 230959
rect 22389 230897 22699 230931
rect 22389 230869 22437 230897
rect 22465 230869 22499 230897
rect 22527 230869 22561 230897
rect 22589 230869 22623 230897
rect 22651 230869 22699 230897
rect 22389 230835 22699 230869
rect 22389 230807 22437 230835
rect 22465 230807 22499 230835
rect 22527 230807 22561 230835
rect 22589 230807 22623 230835
rect 22651 230807 22699 230835
rect 22389 230773 22699 230807
rect 22389 230745 22437 230773
rect 22465 230745 22499 230773
rect 22527 230745 22561 230773
rect 22589 230745 22623 230773
rect 22651 230745 22699 230773
rect 22389 221959 22699 230745
rect 24904 230959 25064 230976
rect 24904 230931 24939 230959
rect 24967 230931 25001 230959
rect 25029 230931 25064 230959
rect 24904 230897 25064 230931
rect 24904 230869 24939 230897
rect 24967 230869 25001 230897
rect 25029 230869 25064 230897
rect 24904 230835 25064 230869
rect 24904 230807 24939 230835
rect 24967 230807 25001 230835
rect 25029 230807 25064 230835
rect 24904 230773 25064 230807
rect 24904 230745 24939 230773
rect 24967 230745 25001 230773
rect 25029 230745 25064 230773
rect 24904 230728 25064 230745
rect 29529 227959 29839 236745
rect 29529 227931 29577 227959
rect 29605 227931 29639 227959
rect 29667 227931 29701 227959
rect 29729 227931 29763 227959
rect 29791 227931 29839 227959
rect 29529 227897 29839 227931
rect 29529 227869 29577 227897
rect 29605 227869 29639 227897
rect 29667 227869 29701 227897
rect 29729 227869 29763 227897
rect 29791 227869 29839 227897
rect 29529 227835 29839 227869
rect 29529 227807 29577 227835
rect 29605 227807 29639 227835
rect 29667 227807 29701 227835
rect 29729 227807 29763 227835
rect 29791 227807 29839 227835
rect 29529 227773 29839 227807
rect 29529 227745 29577 227773
rect 29605 227745 29639 227773
rect 29667 227745 29701 227773
rect 29729 227745 29763 227773
rect 29791 227745 29839 227773
rect 22389 221931 22437 221959
rect 22465 221931 22499 221959
rect 22527 221931 22561 221959
rect 22589 221931 22623 221959
rect 22651 221931 22699 221959
rect 22389 221897 22699 221931
rect 22389 221869 22437 221897
rect 22465 221869 22499 221897
rect 22527 221869 22561 221897
rect 22589 221869 22623 221897
rect 22651 221869 22699 221897
rect 22389 221835 22699 221869
rect 22389 221807 22437 221835
rect 22465 221807 22499 221835
rect 22527 221807 22561 221835
rect 22589 221807 22623 221835
rect 22651 221807 22699 221835
rect 22389 221773 22699 221807
rect 22389 221745 22437 221773
rect 22465 221745 22499 221773
rect 22527 221745 22561 221773
rect 22589 221745 22623 221773
rect 22651 221745 22699 221773
rect 22389 212959 22699 221745
rect 24904 221959 25064 221976
rect 24904 221931 24939 221959
rect 24967 221931 25001 221959
rect 25029 221931 25064 221959
rect 24904 221897 25064 221931
rect 24904 221869 24939 221897
rect 24967 221869 25001 221897
rect 25029 221869 25064 221897
rect 24904 221835 25064 221869
rect 24904 221807 24939 221835
rect 24967 221807 25001 221835
rect 25029 221807 25064 221835
rect 24904 221773 25064 221807
rect 24904 221745 24939 221773
rect 24967 221745 25001 221773
rect 25029 221745 25064 221773
rect 24904 221728 25064 221745
rect 29529 218959 29839 227745
rect 29529 218931 29577 218959
rect 29605 218931 29639 218959
rect 29667 218931 29701 218959
rect 29729 218931 29763 218959
rect 29791 218931 29839 218959
rect 29529 218897 29839 218931
rect 29529 218869 29577 218897
rect 29605 218869 29639 218897
rect 29667 218869 29701 218897
rect 29729 218869 29763 218897
rect 29791 218869 29839 218897
rect 29529 218835 29839 218869
rect 29529 218807 29577 218835
rect 29605 218807 29639 218835
rect 29667 218807 29701 218835
rect 29729 218807 29763 218835
rect 29791 218807 29839 218835
rect 29529 218773 29839 218807
rect 29529 218745 29577 218773
rect 29605 218745 29639 218773
rect 29667 218745 29701 218773
rect 29729 218745 29763 218773
rect 29791 218745 29839 218773
rect 22389 212931 22437 212959
rect 22465 212931 22499 212959
rect 22527 212931 22561 212959
rect 22589 212931 22623 212959
rect 22651 212931 22699 212959
rect 22389 212897 22699 212931
rect 22389 212869 22437 212897
rect 22465 212869 22499 212897
rect 22527 212869 22561 212897
rect 22589 212869 22623 212897
rect 22651 212869 22699 212897
rect 22389 212835 22699 212869
rect 22389 212807 22437 212835
rect 22465 212807 22499 212835
rect 22527 212807 22561 212835
rect 22589 212807 22623 212835
rect 22651 212807 22699 212835
rect 22389 212773 22699 212807
rect 22389 212745 22437 212773
rect 22465 212745 22499 212773
rect 22527 212745 22561 212773
rect 22589 212745 22623 212773
rect 22651 212745 22699 212773
rect 22389 203959 22699 212745
rect 24904 212959 25064 212976
rect 24904 212931 24939 212959
rect 24967 212931 25001 212959
rect 25029 212931 25064 212959
rect 24904 212897 25064 212931
rect 24904 212869 24939 212897
rect 24967 212869 25001 212897
rect 25029 212869 25064 212897
rect 24904 212835 25064 212869
rect 24904 212807 24939 212835
rect 24967 212807 25001 212835
rect 25029 212807 25064 212835
rect 24904 212773 25064 212807
rect 24904 212745 24939 212773
rect 24967 212745 25001 212773
rect 25029 212745 25064 212773
rect 24904 212728 25064 212745
rect 29529 209959 29839 218745
rect 29529 209931 29577 209959
rect 29605 209931 29639 209959
rect 29667 209931 29701 209959
rect 29729 209931 29763 209959
rect 29791 209931 29839 209959
rect 29529 209897 29839 209931
rect 29529 209869 29577 209897
rect 29605 209869 29639 209897
rect 29667 209869 29701 209897
rect 29729 209869 29763 209897
rect 29791 209869 29839 209897
rect 29529 209835 29839 209869
rect 29529 209807 29577 209835
rect 29605 209807 29639 209835
rect 29667 209807 29701 209835
rect 29729 209807 29763 209835
rect 29791 209807 29839 209835
rect 29529 209773 29839 209807
rect 29529 209745 29577 209773
rect 29605 209745 29639 209773
rect 29667 209745 29701 209773
rect 29729 209745 29763 209773
rect 29791 209745 29839 209773
rect 22389 203931 22437 203959
rect 22465 203931 22499 203959
rect 22527 203931 22561 203959
rect 22589 203931 22623 203959
rect 22651 203931 22699 203959
rect 22389 203897 22699 203931
rect 22389 203869 22437 203897
rect 22465 203869 22499 203897
rect 22527 203869 22561 203897
rect 22589 203869 22623 203897
rect 22651 203869 22699 203897
rect 22389 203835 22699 203869
rect 22389 203807 22437 203835
rect 22465 203807 22499 203835
rect 22527 203807 22561 203835
rect 22589 203807 22623 203835
rect 22651 203807 22699 203835
rect 22389 203773 22699 203807
rect 22389 203745 22437 203773
rect 22465 203745 22499 203773
rect 22527 203745 22561 203773
rect 22589 203745 22623 203773
rect 22651 203745 22699 203773
rect 22389 194959 22699 203745
rect 24904 203959 25064 203976
rect 24904 203931 24939 203959
rect 24967 203931 25001 203959
rect 25029 203931 25064 203959
rect 24904 203897 25064 203931
rect 24904 203869 24939 203897
rect 24967 203869 25001 203897
rect 25029 203869 25064 203897
rect 24904 203835 25064 203869
rect 24904 203807 24939 203835
rect 24967 203807 25001 203835
rect 25029 203807 25064 203835
rect 24904 203773 25064 203807
rect 24904 203745 24939 203773
rect 24967 203745 25001 203773
rect 25029 203745 25064 203773
rect 24904 203728 25064 203745
rect 29529 200959 29839 209745
rect 29529 200931 29577 200959
rect 29605 200931 29639 200959
rect 29667 200931 29701 200959
rect 29729 200931 29763 200959
rect 29791 200931 29839 200959
rect 29529 200897 29839 200931
rect 29529 200869 29577 200897
rect 29605 200869 29639 200897
rect 29667 200869 29701 200897
rect 29729 200869 29763 200897
rect 29791 200869 29839 200897
rect 29529 200835 29839 200869
rect 29529 200807 29577 200835
rect 29605 200807 29639 200835
rect 29667 200807 29701 200835
rect 29729 200807 29763 200835
rect 29791 200807 29839 200835
rect 29529 200773 29839 200807
rect 29529 200745 29577 200773
rect 29605 200745 29639 200773
rect 29667 200745 29701 200773
rect 29729 200745 29763 200773
rect 29791 200745 29839 200773
rect 22389 194931 22437 194959
rect 22465 194931 22499 194959
rect 22527 194931 22561 194959
rect 22589 194931 22623 194959
rect 22651 194931 22699 194959
rect 22389 194897 22699 194931
rect 22389 194869 22437 194897
rect 22465 194869 22499 194897
rect 22527 194869 22561 194897
rect 22589 194869 22623 194897
rect 22651 194869 22699 194897
rect 22389 194835 22699 194869
rect 22389 194807 22437 194835
rect 22465 194807 22499 194835
rect 22527 194807 22561 194835
rect 22589 194807 22623 194835
rect 22651 194807 22699 194835
rect 22389 194773 22699 194807
rect 22389 194745 22437 194773
rect 22465 194745 22499 194773
rect 22527 194745 22561 194773
rect 22589 194745 22623 194773
rect 22651 194745 22699 194773
rect 22389 185959 22699 194745
rect 24904 194959 25064 194976
rect 24904 194931 24939 194959
rect 24967 194931 25001 194959
rect 25029 194931 25064 194959
rect 24904 194897 25064 194931
rect 24904 194869 24939 194897
rect 24967 194869 25001 194897
rect 25029 194869 25064 194897
rect 24904 194835 25064 194869
rect 24904 194807 24939 194835
rect 24967 194807 25001 194835
rect 25029 194807 25064 194835
rect 24904 194773 25064 194807
rect 24904 194745 24939 194773
rect 24967 194745 25001 194773
rect 25029 194745 25064 194773
rect 24904 194728 25064 194745
rect 29529 191959 29839 200745
rect 29529 191931 29577 191959
rect 29605 191931 29639 191959
rect 29667 191931 29701 191959
rect 29729 191931 29763 191959
rect 29791 191931 29839 191959
rect 29529 191897 29839 191931
rect 29529 191869 29577 191897
rect 29605 191869 29639 191897
rect 29667 191869 29701 191897
rect 29729 191869 29763 191897
rect 29791 191869 29839 191897
rect 29529 191835 29839 191869
rect 29529 191807 29577 191835
rect 29605 191807 29639 191835
rect 29667 191807 29701 191835
rect 29729 191807 29763 191835
rect 29791 191807 29839 191835
rect 29529 191773 29839 191807
rect 29529 191745 29577 191773
rect 29605 191745 29639 191773
rect 29667 191745 29701 191773
rect 29729 191745 29763 191773
rect 29791 191745 29839 191773
rect 22389 185931 22437 185959
rect 22465 185931 22499 185959
rect 22527 185931 22561 185959
rect 22589 185931 22623 185959
rect 22651 185931 22699 185959
rect 22389 185897 22699 185931
rect 22389 185869 22437 185897
rect 22465 185869 22499 185897
rect 22527 185869 22561 185897
rect 22589 185869 22623 185897
rect 22651 185869 22699 185897
rect 22389 185835 22699 185869
rect 22389 185807 22437 185835
rect 22465 185807 22499 185835
rect 22527 185807 22561 185835
rect 22589 185807 22623 185835
rect 22651 185807 22699 185835
rect 22389 185773 22699 185807
rect 22389 185745 22437 185773
rect 22465 185745 22499 185773
rect 22527 185745 22561 185773
rect 22589 185745 22623 185773
rect 22651 185745 22699 185773
rect 22389 176959 22699 185745
rect 24904 185959 25064 185976
rect 24904 185931 24939 185959
rect 24967 185931 25001 185959
rect 25029 185931 25064 185959
rect 24904 185897 25064 185931
rect 24904 185869 24939 185897
rect 24967 185869 25001 185897
rect 25029 185869 25064 185897
rect 24904 185835 25064 185869
rect 24904 185807 24939 185835
rect 24967 185807 25001 185835
rect 25029 185807 25064 185835
rect 24904 185773 25064 185807
rect 24904 185745 24939 185773
rect 24967 185745 25001 185773
rect 25029 185745 25064 185773
rect 24904 185728 25064 185745
rect 29529 182959 29839 191745
rect 29529 182931 29577 182959
rect 29605 182931 29639 182959
rect 29667 182931 29701 182959
rect 29729 182931 29763 182959
rect 29791 182931 29839 182959
rect 29529 182897 29839 182931
rect 29529 182869 29577 182897
rect 29605 182869 29639 182897
rect 29667 182869 29701 182897
rect 29729 182869 29763 182897
rect 29791 182869 29839 182897
rect 29529 182835 29839 182869
rect 29529 182807 29577 182835
rect 29605 182807 29639 182835
rect 29667 182807 29701 182835
rect 29729 182807 29763 182835
rect 29791 182807 29839 182835
rect 29529 182773 29839 182807
rect 29529 182745 29577 182773
rect 29605 182745 29639 182773
rect 29667 182745 29701 182773
rect 29729 182745 29763 182773
rect 29791 182745 29839 182773
rect 22389 176931 22437 176959
rect 22465 176931 22499 176959
rect 22527 176931 22561 176959
rect 22589 176931 22623 176959
rect 22651 176931 22699 176959
rect 22389 176897 22699 176931
rect 22389 176869 22437 176897
rect 22465 176869 22499 176897
rect 22527 176869 22561 176897
rect 22589 176869 22623 176897
rect 22651 176869 22699 176897
rect 22389 176835 22699 176869
rect 22389 176807 22437 176835
rect 22465 176807 22499 176835
rect 22527 176807 22561 176835
rect 22589 176807 22623 176835
rect 22651 176807 22699 176835
rect 22389 176773 22699 176807
rect 22389 176745 22437 176773
rect 22465 176745 22499 176773
rect 22527 176745 22561 176773
rect 22589 176745 22623 176773
rect 22651 176745 22699 176773
rect 22389 167959 22699 176745
rect 24904 176959 25064 176976
rect 24904 176931 24939 176959
rect 24967 176931 25001 176959
rect 25029 176931 25064 176959
rect 24904 176897 25064 176931
rect 24904 176869 24939 176897
rect 24967 176869 25001 176897
rect 25029 176869 25064 176897
rect 24904 176835 25064 176869
rect 24904 176807 24939 176835
rect 24967 176807 25001 176835
rect 25029 176807 25064 176835
rect 24904 176773 25064 176807
rect 24904 176745 24939 176773
rect 24967 176745 25001 176773
rect 25029 176745 25064 176773
rect 24904 176728 25064 176745
rect 29529 173959 29839 182745
rect 29529 173931 29577 173959
rect 29605 173931 29639 173959
rect 29667 173931 29701 173959
rect 29729 173931 29763 173959
rect 29791 173931 29839 173959
rect 29529 173897 29839 173931
rect 29529 173869 29577 173897
rect 29605 173869 29639 173897
rect 29667 173869 29701 173897
rect 29729 173869 29763 173897
rect 29791 173869 29839 173897
rect 29529 173835 29839 173869
rect 29529 173807 29577 173835
rect 29605 173807 29639 173835
rect 29667 173807 29701 173835
rect 29729 173807 29763 173835
rect 29791 173807 29839 173835
rect 29529 173773 29839 173807
rect 29529 173745 29577 173773
rect 29605 173745 29639 173773
rect 29667 173745 29701 173773
rect 29729 173745 29763 173773
rect 29791 173745 29839 173773
rect 22389 167931 22437 167959
rect 22465 167931 22499 167959
rect 22527 167931 22561 167959
rect 22589 167931 22623 167959
rect 22651 167931 22699 167959
rect 22389 167897 22699 167931
rect 22389 167869 22437 167897
rect 22465 167869 22499 167897
rect 22527 167869 22561 167897
rect 22589 167869 22623 167897
rect 22651 167869 22699 167897
rect 22389 167835 22699 167869
rect 22389 167807 22437 167835
rect 22465 167807 22499 167835
rect 22527 167807 22561 167835
rect 22589 167807 22623 167835
rect 22651 167807 22699 167835
rect 22389 167773 22699 167807
rect 22389 167745 22437 167773
rect 22465 167745 22499 167773
rect 22527 167745 22561 167773
rect 22589 167745 22623 167773
rect 22651 167745 22699 167773
rect 22389 158959 22699 167745
rect 24904 167959 25064 167976
rect 24904 167931 24939 167959
rect 24967 167931 25001 167959
rect 25029 167931 25064 167959
rect 24904 167897 25064 167931
rect 24904 167869 24939 167897
rect 24967 167869 25001 167897
rect 25029 167869 25064 167897
rect 24904 167835 25064 167869
rect 24904 167807 24939 167835
rect 24967 167807 25001 167835
rect 25029 167807 25064 167835
rect 24904 167773 25064 167807
rect 24904 167745 24939 167773
rect 24967 167745 25001 167773
rect 25029 167745 25064 167773
rect 24904 167728 25064 167745
rect 29529 164959 29839 173745
rect 29529 164931 29577 164959
rect 29605 164931 29639 164959
rect 29667 164931 29701 164959
rect 29729 164931 29763 164959
rect 29791 164931 29839 164959
rect 29529 164897 29839 164931
rect 29529 164869 29577 164897
rect 29605 164869 29639 164897
rect 29667 164869 29701 164897
rect 29729 164869 29763 164897
rect 29791 164869 29839 164897
rect 29529 164835 29839 164869
rect 29529 164807 29577 164835
rect 29605 164807 29639 164835
rect 29667 164807 29701 164835
rect 29729 164807 29763 164835
rect 29791 164807 29839 164835
rect 29529 164773 29839 164807
rect 29529 164745 29577 164773
rect 29605 164745 29639 164773
rect 29667 164745 29701 164773
rect 29729 164745 29763 164773
rect 29791 164745 29839 164773
rect 22389 158931 22437 158959
rect 22465 158931 22499 158959
rect 22527 158931 22561 158959
rect 22589 158931 22623 158959
rect 22651 158931 22699 158959
rect 22389 158897 22699 158931
rect 22389 158869 22437 158897
rect 22465 158869 22499 158897
rect 22527 158869 22561 158897
rect 22589 158869 22623 158897
rect 22651 158869 22699 158897
rect 22389 158835 22699 158869
rect 22389 158807 22437 158835
rect 22465 158807 22499 158835
rect 22527 158807 22561 158835
rect 22589 158807 22623 158835
rect 22651 158807 22699 158835
rect 22389 158773 22699 158807
rect 22389 158745 22437 158773
rect 22465 158745 22499 158773
rect 22527 158745 22561 158773
rect 22589 158745 22623 158773
rect 22651 158745 22699 158773
rect 22389 149959 22699 158745
rect 24904 158959 25064 158976
rect 24904 158931 24939 158959
rect 24967 158931 25001 158959
rect 25029 158931 25064 158959
rect 24904 158897 25064 158931
rect 24904 158869 24939 158897
rect 24967 158869 25001 158897
rect 25029 158869 25064 158897
rect 24904 158835 25064 158869
rect 24904 158807 24939 158835
rect 24967 158807 25001 158835
rect 25029 158807 25064 158835
rect 24904 158773 25064 158807
rect 24904 158745 24939 158773
rect 24967 158745 25001 158773
rect 25029 158745 25064 158773
rect 24904 158728 25064 158745
rect 29529 155959 29839 164745
rect 29529 155931 29577 155959
rect 29605 155931 29639 155959
rect 29667 155931 29701 155959
rect 29729 155931 29763 155959
rect 29791 155931 29839 155959
rect 29529 155897 29839 155931
rect 29529 155869 29577 155897
rect 29605 155869 29639 155897
rect 29667 155869 29701 155897
rect 29729 155869 29763 155897
rect 29791 155869 29839 155897
rect 29529 155835 29839 155869
rect 29529 155807 29577 155835
rect 29605 155807 29639 155835
rect 29667 155807 29701 155835
rect 29729 155807 29763 155835
rect 29791 155807 29839 155835
rect 29529 155773 29839 155807
rect 29529 155745 29577 155773
rect 29605 155745 29639 155773
rect 29667 155745 29701 155773
rect 29729 155745 29763 155773
rect 29791 155745 29839 155773
rect 22389 149931 22437 149959
rect 22465 149931 22499 149959
rect 22527 149931 22561 149959
rect 22589 149931 22623 149959
rect 22651 149931 22699 149959
rect 22389 149897 22699 149931
rect 22389 149869 22437 149897
rect 22465 149869 22499 149897
rect 22527 149869 22561 149897
rect 22589 149869 22623 149897
rect 22651 149869 22699 149897
rect 22389 149835 22699 149869
rect 22389 149807 22437 149835
rect 22465 149807 22499 149835
rect 22527 149807 22561 149835
rect 22589 149807 22623 149835
rect 22651 149807 22699 149835
rect 22389 149773 22699 149807
rect 22389 149745 22437 149773
rect 22465 149745 22499 149773
rect 22527 149745 22561 149773
rect 22589 149745 22623 149773
rect 22651 149745 22699 149773
rect 22389 140959 22699 149745
rect 24904 149959 25064 149976
rect 24904 149931 24939 149959
rect 24967 149931 25001 149959
rect 25029 149931 25064 149959
rect 24904 149897 25064 149931
rect 24904 149869 24939 149897
rect 24967 149869 25001 149897
rect 25029 149869 25064 149897
rect 24904 149835 25064 149869
rect 24904 149807 24939 149835
rect 24967 149807 25001 149835
rect 25029 149807 25064 149835
rect 24904 149773 25064 149807
rect 24904 149745 24939 149773
rect 24967 149745 25001 149773
rect 25029 149745 25064 149773
rect 24904 149728 25064 149745
rect 29529 146959 29839 155745
rect 29529 146931 29577 146959
rect 29605 146931 29639 146959
rect 29667 146931 29701 146959
rect 29729 146931 29763 146959
rect 29791 146931 29839 146959
rect 29529 146897 29839 146931
rect 29529 146869 29577 146897
rect 29605 146869 29639 146897
rect 29667 146869 29701 146897
rect 29729 146869 29763 146897
rect 29791 146869 29839 146897
rect 29529 146835 29839 146869
rect 29529 146807 29577 146835
rect 29605 146807 29639 146835
rect 29667 146807 29701 146835
rect 29729 146807 29763 146835
rect 29791 146807 29839 146835
rect 29529 146773 29839 146807
rect 29529 146745 29577 146773
rect 29605 146745 29639 146773
rect 29667 146745 29701 146773
rect 29729 146745 29763 146773
rect 29791 146745 29839 146773
rect 22389 140931 22437 140959
rect 22465 140931 22499 140959
rect 22527 140931 22561 140959
rect 22589 140931 22623 140959
rect 22651 140931 22699 140959
rect 22389 140897 22699 140931
rect 22389 140869 22437 140897
rect 22465 140869 22499 140897
rect 22527 140869 22561 140897
rect 22589 140869 22623 140897
rect 22651 140869 22699 140897
rect 22389 140835 22699 140869
rect 22389 140807 22437 140835
rect 22465 140807 22499 140835
rect 22527 140807 22561 140835
rect 22589 140807 22623 140835
rect 22651 140807 22699 140835
rect 22389 140773 22699 140807
rect 22389 140745 22437 140773
rect 22465 140745 22499 140773
rect 22527 140745 22561 140773
rect 22589 140745 22623 140773
rect 22651 140745 22699 140773
rect 22389 131959 22699 140745
rect 24904 140959 25064 140976
rect 24904 140931 24939 140959
rect 24967 140931 25001 140959
rect 25029 140931 25064 140959
rect 24904 140897 25064 140931
rect 24904 140869 24939 140897
rect 24967 140869 25001 140897
rect 25029 140869 25064 140897
rect 24904 140835 25064 140869
rect 24904 140807 24939 140835
rect 24967 140807 25001 140835
rect 25029 140807 25064 140835
rect 24904 140773 25064 140807
rect 24904 140745 24939 140773
rect 24967 140745 25001 140773
rect 25029 140745 25064 140773
rect 24904 140728 25064 140745
rect 29529 137959 29839 146745
rect 29529 137931 29577 137959
rect 29605 137931 29639 137959
rect 29667 137931 29701 137959
rect 29729 137931 29763 137959
rect 29791 137931 29839 137959
rect 29529 137897 29839 137931
rect 29529 137869 29577 137897
rect 29605 137869 29639 137897
rect 29667 137869 29701 137897
rect 29729 137869 29763 137897
rect 29791 137869 29839 137897
rect 29529 137835 29839 137869
rect 29529 137807 29577 137835
rect 29605 137807 29639 137835
rect 29667 137807 29701 137835
rect 29729 137807 29763 137835
rect 29791 137807 29839 137835
rect 29529 137773 29839 137807
rect 29529 137745 29577 137773
rect 29605 137745 29639 137773
rect 29667 137745 29701 137773
rect 29729 137745 29763 137773
rect 29791 137745 29839 137773
rect 22389 131931 22437 131959
rect 22465 131931 22499 131959
rect 22527 131931 22561 131959
rect 22589 131931 22623 131959
rect 22651 131931 22699 131959
rect 22389 131897 22699 131931
rect 22389 131869 22437 131897
rect 22465 131869 22499 131897
rect 22527 131869 22561 131897
rect 22589 131869 22623 131897
rect 22651 131869 22699 131897
rect 22389 131835 22699 131869
rect 22389 131807 22437 131835
rect 22465 131807 22499 131835
rect 22527 131807 22561 131835
rect 22589 131807 22623 131835
rect 22651 131807 22699 131835
rect 22389 131773 22699 131807
rect 22389 131745 22437 131773
rect 22465 131745 22499 131773
rect 22527 131745 22561 131773
rect 22589 131745 22623 131773
rect 22651 131745 22699 131773
rect 22389 122959 22699 131745
rect 24904 131959 25064 131976
rect 24904 131931 24939 131959
rect 24967 131931 25001 131959
rect 25029 131931 25064 131959
rect 24904 131897 25064 131931
rect 24904 131869 24939 131897
rect 24967 131869 25001 131897
rect 25029 131869 25064 131897
rect 24904 131835 25064 131869
rect 24904 131807 24939 131835
rect 24967 131807 25001 131835
rect 25029 131807 25064 131835
rect 24904 131773 25064 131807
rect 24904 131745 24939 131773
rect 24967 131745 25001 131773
rect 25029 131745 25064 131773
rect 24904 131728 25064 131745
rect 29529 128959 29839 137745
rect 29529 128931 29577 128959
rect 29605 128931 29639 128959
rect 29667 128931 29701 128959
rect 29729 128931 29763 128959
rect 29791 128931 29839 128959
rect 29529 128897 29839 128931
rect 29529 128869 29577 128897
rect 29605 128869 29639 128897
rect 29667 128869 29701 128897
rect 29729 128869 29763 128897
rect 29791 128869 29839 128897
rect 29529 128835 29839 128869
rect 29529 128807 29577 128835
rect 29605 128807 29639 128835
rect 29667 128807 29701 128835
rect 29729 128807 29763 128835
rect 29791 128807 29839 128835
rect 29529 128773 29839 128807
rect 29529 128745 29577 128773
rect 29605 128745 29639 128773
rect 29667 128745 29701 128773
rect 29729 128745 29763 128773
rect 29791 128745 29839 128773
rect 22389 122931 22437 122959
rect 22465 122931 22499 122959
rect 22527 122931 22561 122959
rect 22589 122931 22623 122959
rect 22651 122931 22699 122959
rect 22389 122897 22699 122931
rect 22389 122869 22437 122897
rect 22465 122869 22499 122897
rect 22527 122869 22561 122897
rect 22589 122869 22623 122897
rect 22651 122869 22699 122897
rect 22389 122835 22699 122869
rect 22389 122807 22437 122835
rect 22465 122807 22499 122835
rect 22527 122807 22561 122835
rect 22589 122807 22623 122835
rect 22651 122807 22699 122835
rect 22389 122773 22699 122807
rect 22389 122745 22437 122773
rect 22465 122745 22499 122773
rect 22527 122745 22561 122773
rect 22589 122745 22623 122773
rect 22651 122745 22699 122773
rect 22389 113959 22699 122745
rect 24904 122959 25064 122976
rect 24904 122931 24939 122959
rect 24967 122931 25001 122959
rect 25029 122931 25064 122959
rect 24904 122897 25064 122931
rect 24904 122869 24939 122897
rect 24967 122869 25001 122897
rect 25029 122869 25064 122897
rect 24904 122835 25064 122869
rect 24904 122807 24939 122835
rect 24967 122807 25001 122835
rect 25029 122807 25064 122835
rect 24904 122773 25064 122807
rect 24904 122745 24939 122773
rect 24967 122745 25001 122773
rect 25029 122745 25064 122773
rect 24904 122728 25064 122745
rect 29529 119959 29839 128745
rect 29529 119931 29577 119959
rect 29605 119931 29639 119959
rect 29667 119931 29701 119959
rect 29729 119931 29763 119959
rect 29791 119931 29839 119959
rect 29529 119897 29839 119931
rect 29529 119869 29577 119897
rect 29605 119869 29639 119897
rect 29667 119869 29701 119897
rect 29729 119869 29763 119897
rect 29791 119869 29839 119897
rect 29529 119835 29839 119869
rect 29529 119807 29577 119835
rect 29605 119807 29639 119835
rect 29667 119807 29701 119835
rect 29729 119807 29763 119835
rect 29791 119807 29839 119835
rect 29529 119773 29839 119807
rect 29529 119745 29577 119773
rect 29605 119745 29639 119773
rect 29667 119745 29701 119773
rect 29729 119745 29763 119773
rect 29791 119745 29839 119773
rect 22389 113931 22437 113959
rect 22465 113931 22499 113959
rect 22527 113931 22561 113959
rect 22589 113931 22623 113959
rect 22651 113931 22699 113959
rect 22389 113897 22699 113931
rect 22389 113869 22437 113897
rect 22465 113869 22499 113897
rect 22527 113869 22561 113897
rect 22589 113869 22623 113897
rect 22651 113869 22699 113897
rect 22389 113835 22699 113869
rect 22389 113807 22437 113835
rect 22465 113807 22499 113835
rect 22527 113807 22561 113835
rect 22589 113807 22623 113835
rect 22651 113807 22699 113835
rect 22389 113773 22699 113807
rect 22389 113745 22437 113773
rect 22465 113745 22499 113773
rect 22527 113745 22561 113773
rect 22589 113745 22623 113773
rect 22651 113745 22699 113773
rect 22389 104959 22699 113745
rect 24904 113959 25064 113976
rect 24904 113931 24939 113959
rect 24967 113931 25001 113959
rect 25029 113931 25064 113959
rect 24904 113897 25064 113931
rect 24904 113869 24939 113897
rect 24967 113869 25001 113897
rect 25029 113869 25064 113897
rect 24904 113835 25064 113869
rect 24904 113807 24939 113835
rect 24967 113807 25001 113835
rect 25029 113807 25064 113835
rect 24904 113773 25064 113807
rect 24904 113745 24939 113773
rect 24967 113745 25001 113773
rect 25029 113745 25064 113773
rect 24904 113728 25064 113745
rect 29529 110959 29839 119745
rect 29529 110931 29577 110959
rect 29605 110931 29639 110959
rect 29667 110931 29701 110959
rect 29729 110931 29763 110959
rect 29791 110931 29839 110959
rect 29529 110897 29839 110931
rect 29529 110869 29577 110897
rect 29605 110869 29639 110897
rect 29667 110869 29701 110897
rect 29729 110869 29763 110897
rect 29791 110869 29839 110897
rect 29529 110835 29839 110869
rect 29529 110807 29577 110835
rect 29605 110807 29639 110835
rect 29667 110807 29701 110835
rect 29729 110807 29763 110835
rect 29791 110807 29839 110835
rect 29529 110773 29839 110807
rect 29529 110745 29577 110773
rect 29605 110745 29639 110773
rect 29667 110745 29701 110773
rect 29729 110745 29763 110773
rect 29791 110745 29839 110773
rect 22389 104931 22437 104959
rect 22465 104931 22499 104959
rect 22527 104931 22561 104959
rect 22589 104931 22623 104959
rect 22651 104931 22699 104959
rect 22389 104897 22699 104931
rect 22389 104869 22437 104897
rect 22465 104869 22499 104897
rect 22527 104869 22561 104897
rect 22589 104869 22623 104897
rect 22651 104869 22699 104897
rect 22389 104835 22699 104869
rect 22389 104807 22437 104835
rect 22465 104807 22499 104835
rect 22527 104807 22561 104835
rect 22589 104807 22623 104835
rect 22651 104807 22699 104835
rect 22389 104773 22699 104807
rect 22389 104745 22437 104773
rect 22465 104745 22499 104773
rect 22527 104745 22561 104773
rect 22589 104745 22623 104773
rect 22651 104745 22699 104773
rect 22389 95959 22699 104745
rect 24904 104959 25064 104976
rect 24904 104931 24939 104959
rect 24967 104931 25001 104959
rect 25029 104931 25064 104959
rect 24904 104897 25064 104931
rect 24904 104869 24939 104897
rect 24967 104869 25001 104897
rect 25029 104869 25064 104897
rect 24904 104835 25064 104869
rect 24904 104807 24939 104835
rect 24967 104807 25001 104835
rect 25029 104807 25064 104835
rect 24904 104773 25064 104807
rect 24904 104745 24939 104773
rect 24967 104745 25001 104773
rect 25029 104745 25064 104773
rect 24904 104728 25064 104745
rect 29529 101959 29839 110745
rect 29529 101931 29577 101959
rect 29605 101931 29639 101959
rect 29667 101931 29701 101959
rect 29729 101931 29763 101959
rect 29791 101931 29839 101959
rect 29529 101897 29839 101931
rect 29529 101869 29577 101897
rect 29605 101869 29639 101897
rect 29667 101869 29701 101897
rect 29729 101869 29763 101897
rect 29791 101869 29839 101897
rect 29529 101835 29839 101869
rect 29529 101807 29577 101835
rect 29605 101807 29639 101835
rect 29667 101807 29701 101835
rect 29729 101807 29763 101835
rect 29791 101807 29839 101835
rect 29529 101773 29839 101807
rect 29529 101745 29577 101773
rect 29605 101745 29639 101773
rect 29667 101745 29701 101773
rect 29729 101745 29763 101773
rect 29791 101745 29839 101773
rect 22389 95931 22437 95959
rect 22465 95931 22499 95959
rect 22527 95931 22561 95959
rect 22589 95931 22623 95959
rect 22651 95931 22699 95959
rect 22389 95897 22699 95931
rect 22389 95869 22437 95897
rect 22465 95869 22499 95897
rect 22527 95869 22561 95897
rect 22589 95869 22623 95897
rect 22651 95869 22699 95897
rect 22389 95835 22699 95869
rect 22389 95807 22437 95835
rect 22465 95807 22499 95835
rect 22527 95807 22561 95835
rect 22589 95807 22623 95835
rect 22651 95807 22699 95835
rect 22389 95773 22699 95807
rect 22389 95745 22437 95773
rect 22465 95745 22499 95773
rect 22527 95745 22561 95773
rect 22589 95745 22623 95773
rect 22651 95745 22699 95773
rect 22389 86959 22699 95745
rect 24904 95959 25064 95976
rect 24904 95931 24939 95959
rect 24967 95931 25001 95959
rect 25029 95931 25064 95959
rect 24904 95897 25064 95931
rect 24904 95869 24939 95897
rect 24967 95869 25001 95897
rect 25029 95869 25064 95897
rect 24904 95835 25064 95869
rect 24904 95807 24939 95835
rect 24967 95807 25001 95835
rect 25029 95807 25064 95835
rect 24904 95773 25064 95807
rect 24904 95745 24939 95773
rect 24967 95745 25001 95773
rect 25029 95745 25064 95773
rect 24904 95728 25064 95745
rect 29529 92959 29839 101745
rect 29529 92931 29577 92959
rect 29605 92931 29639 92959
rect 29667 92931 29701 92959
rect 29729 92931 29763 92959
rect 29791 92931 29839 92959
rect 29529 92897 29839 92931
rect 29529 92869 29577 92897
rect 29605 92869 29639 92897
rect 29667 92869 29701 92897
rect 29729 92869 29763 92897
rect 29791 92869 29839 92897
rect 29529 92835 29839 92869
rect 29529 92807 29577 92835
rect 29605 92807 29639 92835
rect 29667 92807 29701 92835
rect 29729 92807 29763 92835
rect 29791 92807 29839 92835
rect 29529 92773 29839 92807
rect 29529 92745 29577 92773
rect 29605 92745 29639 92773
rect 29667 92745 29701 92773
rect 29729 92745 29763 92773
rect 29791 92745 29839 92773
rect 22389 86931 22437 86959
rect 22465 86931 22499 86959
rect 22527 86931 22561 86959
rect 22589 86931 22623 86959
rect 22651 86931 22699 86959
rect 22389 86897 22699 86931
rect 22389 86869 22437 86897
rect 22465 86869 22499 86897
rect 22527 86869 22561 86897
rect 22589 86869 22623 86897
rect 22651 86869 22699 86897
rect 22389 86835 22699 86869
rect 22389 86807 22437 86835
rect 22465 86807 22499 86835
rect 22527 86807 22561 86835
rect 22589 86807 22623 86835
rect 22651 86807 22699 86835
rect 22389 86773 22699 86807
rect 22389 86745 22437 86773
rect 22465 86745 22499 86773
rect 22527 86745 22561 86773
rect 22589 86745 22623 86773
rect 22651 86745 22699 86773
rect 22389 77959 22699 86745
rect 24904 86959 25064 86976
rect 24904 86931 24939 86959
rect 24967 86931 25001 86959
rect 25029 86931 25064 86959
rect 24904 86897 25064 86931
rect 24904 86869 24939 86897
rect 24967 86869 25001 86897
rect 25029 86869 25064 86897
rect 24904 86835 25064 86869
rect 24904 86807 24939 86835
rect 24967 86807 25001 86835
rect 25029 86807 25064 86835
rect 24904 86773 25064 86807
rect 24904 86745 24939 86773
rect 24967 86745 25001 86773
rect 25029 86745 25064 86773
rect 24904 86728 25064 86745
rect 29529 83959 29839 92745
rect 29529 83931 29577 83959
rect 29605 83931 29639 83959
rect 29667 83931 29701 83959
rect 29729 83931 29763 83959
rect 29791 83931 29839 83959
rect 29529 83897 29839 83931
rect 29529 83869 29577 83897
rect 29605 83869 29639 83897
rect 29667 83869 29701 83897
rect 29729 83869 29763 83897
rect 29791 83869 29839 83897
rect 29529 83835 29839 83869
rect 29529 83807 29577 83835
rect 29605 83807 29639 83835
rect 29667 83807 29701 83835
rect 29729 83807 29763 83835
rect 29791 83807 29839 83835
rect 29529 83773 29839 83807
rect 29529 83745 29577 83773
rect 29605 83745 29639 83773
rect 29667 83745 29701 83773
rect 29729 83745 29763 83773
rect 29791 83745 29839 83773
rect 22389 77931 22437 77959
rect 22465 77931 22499 77959
rect 22527 77931 22561 77959
rect 22589 77931 22623 77959
rect 22651 77931 22699 77959
rect 22389 77897 22699 77931
rect 22389 77869 22437 77897
rect 22465 77869 22499 77897
rect 22527 77869 22561 77897
rect 22589 77869 22623 77897
rect 22651 77869 22699 77897
rect 22389 77835 22699 77869
rect 22389 77807 22437 77835
rect 22465 77807 22499 77835
rect 22527 77807 22561 77835
rect 22589 77807 22623 77835
rect 22651 77807 22699 77835
rect 22389 77773 22699 77807
rect 22389 77745 22437 77773
rect 22465 77745 22499 77773
rect 22527 77745 22561 77773
rect 22589 77745 22623 77773
rect 22651 77745 22699 77773
rect 22389 68959 22699 77745
rect 24904 77959 25064 77976
rect 24904 77931 24939 77959
rect 24967 77931 25001 77959
rect 25029 77931 25064 77959
rect 24904 77897 25064 77931
rect 24904 77869 24939 77897
rect 24967 77869 25001 77897
rect 25029 77869 25064 77897
rect 24904 77835 25064 77869
rect 24904 77807 24939 77835
rect 24967 77807 25001 77835
rect 25029 77807 25064 77835
rect 24904 77773 25064 77807
rect 24904 77745 24939 77773
rect 24967 77745 25001 77773
rect 25029 77745 25064 77773
rect 24904 77728 25064 77745
rect 29529 74959 29839 83745
rect 29529 74931 29577 74959
rect 29605 74931 29639 74959
rect 29667 74931 29701 74959
rect 29729 74931 29763 74959
rect 29791 74931 29839 74959
rect 29529 74897 29839 74931
rect 29529 74869 29577 74897
rect 29605 74869 29639 74897
rect 29667 74869 29701 74897
rect 29729 74869 29763 74897
rect 29791 74869 29839 74897
rect 29529 74835 29839 74869
rect 29529 74807 29577 74835
rect 29605 74807 29639 74835
rect 29667 74807 29701 74835
rect 29729 74807 29763 74835
rect 29791 74807 29839 74835
rect 29529 74773 29839 74807
rect 29529 74745 29577 74773
rect 29605 74745 29639 74773
rect 29667 74745 29701 74773
rect 29729 74745 29763 74773
rect 29791 74745 29839 74773
rect 22389 68931 22437 68959
rect 22465 68931 22499 68959
rect 22527 68931 22561 68959
rect 22589 68931 22623 68959
rect 22651 68931 22699 68959
rect 22389 68897 22699 68931
rect 22389 68869 22437 68897
rect 22465 68869 22499 68897
rect 22527 68869 22561 68897
rect 22589 68869 22623 68897
rect 22651 68869 22699 68897
rect 22389 68835 22699 68869
rect 22389 68807 22437 68835
rect 22465 68807 22499 68835
rect 22527 68807 22561 68835
rect 22589 68807 22623 68835
rect 22651 68807 22699 68835
rect 22389 68773 22699 68807
rect 22389 68745 22437 68773
rect 22465 68745 22499 68773
rect 22527 68745 22561 68773
rect 22589 68745 22623 68773
rect 22651 68745 22699 68773
rect 22389 59959 22699 68745
rect 24904 68959 25064 68976
rect 24904 68931 24939 68959
rect 24967 68931 25001 68959
rect 25029 68931 25064 68959
rect 24904 68897 25064 68931
rect 24904 68869 24939 68897
rect 24967 68869 25001 68897
rect 25029 68869 25064 68897
rect 24904 68835 25064 68869
rect 24904 68807 24939 68835
rect 24967 68807 25001 68835
rect 25029 68807 25064 68835
rect 24904 68773 25064 68807
rect 24904 68745 24939 68773
rect 24967 68745 25001 68773
rect 25029 68745 25064 68773
rect 24904 68728 25064 68745
rect 29529 65959 29839 74745
rect 29529 65931 29577 65959
rect 29605 65931 29639 65959
rect 29667 65931 29701 65959
rect 29729 65931 29763 65959
rect 29791 65931 29839 65959
rect 29529 65897 29839 65931
rect 29529 65869 29577 65897
rect 29605 65869 29639 65897
rect 29667 65869 29701 65897
rect 29729 65869 29763 65897
rect 29791 65869 29839 65897
rect 29529 65835 29839 65869
rect 29529 65807 29577 65835
rect 29605 65807 29639 65835
rect 29667 65807 29701 65835
rect 29729 65807 29763 65835
rect 29791 65807 29839 65835
rect 29529 65773 29839 65807
rect 29529 65745 29577 65773
rect 29605 65745 29639 65773
rect 29667 65745 29701 65773
rect 29729 65745 29763 65773
rect 29791 65745 29839 65773
rect 22389 59931 22437 59959
rect 22465 59931 22499 59959
rect 22527 59931 22561 59959
rect 22589 59931 22623 59959
rect 22651 59931 22699 59959
rect 22389 59897 22699 59931
rect 22389 59869 22437 59897
rect 22465 59869 22499 59897
rect 22527 59869 22561 59897
rect 22589 59869 22623 59897
rect 22651 59869 22699 59897
rect 22389 59835 22699 59869
rect 22389 59807 22437 59835
rect 22465 59807 22499 59835
rect 22527 59807 22561 59835
rect 22589 59807 22623 59835
rect 22651 59807 22699 59835
rect 22389 59773 22699 59807
rect 22389 59745 22437 59773
rect 22465 59745 22499 59773
rect 22527 59745 22561 59773
rect 22589 59745 22623 59773
rect 22651 59745 22699 59773
rect 22389 50959 22699 59745
rect 24904 59959 25064 59976
rect 24904 59931 24939 59959
rect 24967 59931 25001 59959
rect 25029 59931 25064 59959
rect 24904 59897 25064 59931
rect 24904 59869 24939 59897
rect 24967 59869 25001 59897
rect 25029 59869 25064 59897
rect 24904 59835 25064 59869
rect 24904 59807 24939 59835
rect 24967 59807 25001 59835
rect 25029 59807 25064 59835
rect 24904 59773 25064 59807
rect 24904 59745 24939 59773
rect 24967 59745 25001 59773
rect 25029 59745 25064 59773
rect 24904 59728 25064 59745
rect 29529 56959 29839 65745
rect 29529 56931 29577 56959
rect 29605 56931 29639 56959
rect 29667 56931 29701 56959
rect 29729 56931 29763 56959
rect 29791 56931 29839 56959
rect 29529 56897 29839 56931
rect 29529 56869 29577 56897
rect 29605 56869 29639 56897
rect 29667 56869 29701 56897
rect 29729 56869 29763 56897
rect 29791 56869 29839 56897
rect 29529 56835 29839 56869
rect 29529 56807 29577 56835
rect 29605 56807 29639 56835
rect 29667 56807 29701 56835
rect 29729 56807 29763 56835
rect 29791 56807 29839 56835
rect 29529 56773 29839 56807
rect 29529 56745 29577 56773
rect 29605 56745 29639 56773
rect 29667 56745 29701 56773
rect 29729 56745 29763 56773
rect 29791 56745 29839 56773
rect 22389 50931 22437 50959
rect 22465 50931 22499 50959
rect 22527 50931 22561 50959
rect 22589 50931 22623 50959
rect 22651 50931 22699 50959
rect 22389 50897 22699 50931
rect 22389 50869 22437 50897
rect 22465 50869 22499 50897
rect 22527 50869 22561 50897
rect 22589 50869 22623 50897
rect 22651 50869 22699 50897
rect 22389 50835 22699 50869
rect 22389 50807 22437 50835
rect 22465 50807 22499 50835
rect 22527 50807 22561 50835
rect 22589 50807 22623 50835
rect 22651 50807 22699 50835
rect 22389 50773 22699 50807
rect 22389 50745 22437 50773
rect 22465 50745 22499 50773
rect 22527 50745 22561 50773
rect 22589 50745 22623 50773
rect 22651 50745 22699 50773
rect 22389 41959 22699 50745
rect 24904 50959 25064 50976
rect 24904 50931 24939 50959
rect 24967 50931 25001 50959
rect 25029 50931 25064 50959
rect 24904 50897 25064 50931
rect 24904 50869 24939 50897
rect 24967 50869 25001 50897
rect 25029 50869 25064 50897
rect 24904 50835 25064 50869
rect 24904 50807 24939 50835
rect 24967 50807 25001 50835
rect 25029 50807 25064 50835
rect 24904 50773 25064 50807
rect 24904 50745 24939 50773
rect 24967 50745 25001 50773
rect 25029 50745 25064 50773
rect 24904 50728 25064 50745
rect 29529 47959 29839 56745
rect 29529 47931 29577 47959
rect 29605 47931 29639 47959
rect 29667 47931 29701 47959
rect 29729 47931 29763 47959
rect 29791 47931 29839 47959
rect 29529 47897 29839 47931
rect 29529 47869 29577 47897
rect 29605 47869 29639 47897
rect 29667 47869 29701 47897
rect 29729 47869 29763 47897
rect 29791 47869 29839 47897
rect 29529 47835 29839 47869
rect 29529 47807 29577 47835
rect 29605 47807 29639 47835
rect 29667 47807 29701 47835
rect 29729 47807 29763 47835
rect 29791 47807 29839 47835
rect 29529 47773 29839 47807
rect 29529 47745 29577 47773
rect 29605 47745 29639 47773
rect 29667 47745 29701 47773
rect 29729 47745 29763 47773
rect 29791 47745 29839 47773
rect 22389 41931 22437 41959
rect 22465 41931 22499 41959
rect 22527 41931 22561 41959
rect 22589 41931 22623 41959
rect 22651 41931 22699 41959
rect 22389 41897 22699 41931
rect 22389 41869 22437 41897
rect 22465 41869 22499 41897
rect 22527 41869 22561 41897
rect 22589 41869 22623 41897
rect 22651 41869 22699 41897
rect 22389 41835 22699 41869
rect 22389 41807 22437 41835
rect 22465 41807 22499 41835
rect 22527 41807 22561 41835
rect 22589 41807 22623 41835
rect 22651 41807 22699 41835
rect 22389 41773 22699 41807
rect 22389 41745 22437 41773
rect 22465 41745 22499 41773
rect 22527 41745 22561 41773
rect 22589 41745 22623 41773
rect 22651 41745 22699 41773
rect 22389 32959 22699 41745
rect 24904 41959 25064 41976
rect 24904 41931 24939 41959
rect 24967 41931 25001 41959
rect 25029 41931 25064 41959
rect 24904 41897 25064 41931
rect 24904 41869 24939 41897
rect 24967 41869 25001 41897
rect 25029 41869 25064 41897
rect 24904 41835 25064 41869
rect 24904 41807 24939 41835
rect 24967 41807 25001 41835
rect 25029 41807 25064 41835
rect 24904 41773 25064 41807
rect 24904 41745 24939 41773
rect 24967 41745 25001 41773
rect 25029 41745 25064 41773
rect 24904 41728 25064 41745
rect 29529 38959 29839 47745
rect 29529 38931 29577 38959
rect 29605 38931 29639 38959
rect 29667 38931 29701 38959
rect 29729 38931 29763 38959
rect 29791 38931 29839 38959
rect 29529 38897 29839 38931
rect 29529 38869 29577 38897
rect 29605 38869 29639 38897
rect 29667 38869 29701 38897
rect 29729 38869 29763 38897
rect 29791 38869 29839 38897
rect 29529 38835 29839 38869
rect 29529 38807 29577 38835
rect 29605 38807 29639 38835
rect 29667 38807 29701 38835
rect 29729 38807 29763 38835
rect 29791 38807 29839 38835
rect 29529 38773 29839 38807
rect 29529 38745 29577 38773
rect 29605 38745 29639 38773
rect 29667 38745 29701 38773
rect 29729 38745 29763 38773
rect 29791 38745 29839 38773
rect 22389 32931 22437 32959
rect 22465 32931 22499 32959
rect 22527 32931 22561 32959
rect 22589 32931 22623 32959
rect 22651 32931 22699 32959
rect 22389 32897 22699 32931
rect 22389 32869 22437 32897
rect 22465 32869 22499 32897
rect 22527 32869 22561 32897
rect 22589 32869 22623 32897
rect 22651 32869 22699 32897
rect 22389 32835 22699 32869
rect 22389 32807 22437 32835
rect 22465 32807 22499 32835
rect 22527 32807 22561 32835
rect 22589 32807 22623 32835
rect 22651 32807 22699 32835
rect 22389 32773 22699 32807
rect 22389 32745 22437 32773
rect 22465 32745 22499 32773
rect 22527 32745 22561 32773
rect 22589 32745 22623 32773
rect 22651 32745 22699 32773
rect 22389 23959 22699 32745
rect 24904 32959 25064 32976
rect 24904 32931 24939 32959
rect 24967 32931 25001 32959
rect 25029 32931 25064 32959
rect 24904 32897 25064 32931
rect 24904 32869 24939 32897
rect 24967 32869 25001 32897
rect 25029 32869 25064 32897
rect 24904 32835 25064 32869
rect 24904 32807 24939 32835
rect 24967 32807 25001 32835
rect 25029 32807 25064 32835
rect 24904 32773 25064 32807
rect 24904 32745 24939 32773
rect 24967 32745 25001 32773
rect 25029 32745 25064 32773
rect 24904 32728 25064 32745
rect 29529 29959 29839 38745
rect 29529 29931 29577 29959
rect 29605 29931 29639 29959
rect 29667 29931 29701 29959
rect 29729 29931 29763 29959
rect 29791 29931 29839 29959
rect 29529 29897 29839 29931
rect 29529 29869 29577 29897
rect 29605 29869 29639 29897
rect 29667 29869 29701 29897
rect 29729 29869 29763 29897
rect 29791 29869 29839 29897
rect 29529 29835 29839 29869
rect 29529 29807 29577 29835
rect 29605 29807 29639 29835
rect 29667 29807 29701 29835
rect 29729 29807 29763 29835
rect 29791 29807 29839 29835
rect 29529 29773 29839 29807
rect 29529 29745 29577 29773
rect 29605 29745 29639 29773
rect 29667 29745 29701 29773
rect 29729 29745 29763 29773
rect 29791 29745 29839 29773
rect 22389 23931 22437 23959
rect 22465 23931 22499 23959
rect 22527 23931 22561 23959
rect 22589 23931 22623 23959
rect 22651 23931 22699 23959
rect 22389 23897 22699 23931
rect 22389 23869 22437 23897
rect 22465 23869 22499 23897
rect 22527 23869 22561 23897
rect 22589 23869 22623 23897
rect 22651 23869 22699 23897
rect 22389 23835 22699 23869
rect 22389 23807 22437 23835
rect 22465 23807 22499 23835
rect 22527 23807 22561 23835
rect 22589 23807 22623 23835
rect 22651 23807 22699 23835
rect 22389 23773 22699 23807
rect 22389 23745 22437 23773
rect 22465 23745 22499 23773
rect 22527 23745 22561 23773
rect 22589 23745 22623 23773
rect 22651 23745 22699 23773
rect 22389 14959 22699 23745
rect 24904 23959 25064 23976
rect 24904 23931 24939 23959
rect 24967 23931 25001 23959
rect 25029 23931 25064 23959
rect 24904 23897 25064 23931
rect 24904 23869 24939 23897
rect 24967 23869 25001 23897
rect 25029 23869 25064 23897
rect 24904 23835 25064 23869
rect 24904 23807 24939 23835
rect 24967 23807 25001 23835
rect 25029 23807 25064 23835
rect 24904 23773 25064 23807
rect 24904 23745 24939 23773
rect 24967 23745 25001 23773
rect 25029 23745 25064 23773
rect 24904 23728 25064 23745
rect 22389 14931 22437 14959
rect 22465 14931 22499 14959
rect 22527 14931 22561 14959
rect 22589 14931 22623 14959
rect 22651 14931 22699 14959
rect 22389 14897 22699 14931
rect 22389 14869 22437 14897
rect 22465 14869 22499 14897
rect 22527 14869 22561 14897
rect 22589 14869 22623 14897
rect 22651 14869 22699 14897
rect 22389 14835 22699 14869
rect 22389 14807 22437 14835
rect 22465 14807 22499 14835
rect 22527 14807 22561 14835
rect 22589 14807 22623 14835
rect 22651 14807 22699 14835
rect 22389 14773 22699 14807
rect 22389 14745 22437 14773
rect 22465 14745 22499 14773
rect 22527 14745 22561 14773
rect 22589 14745 22623 14773
rect 22651 14745 22699 14773
rect 22389 5959 22699 14745
rect 22389 5931 22437 5959
rect 22465 5931 22499 5959
rect 22527 5931 22561 5959
rect 22589 5931 22623 5959
rect 22651 5931 22699 5959
rect 22389 5897 22699 5931
rect 22389 5869 22437 5897
rect 22465 5869 22499 5897
rect 22527 5869 22561 5897
rect 22589 5869 22623 5897
rect 22651 5869 22699 5897
rect 22389 5835 22699 5869
rect 22389 5807 22437 5835
rect 22465 5807 22499 5835
rect 22527 5807 22561 5835
rect 22589 5807 22623 5835
rect 22651 5807 22699 5835
rect 22389 5773 22699 5807
rect 22389 5745 22437 5773
rect 22465 5745 22499 5773
rect 22527 5745 22561 5773
rect 22589 5745 22623 5773
rect 22651 5745 22699 5773
rect 22389 424 22699 5745
rect 22389 396 22437 424
rect 22465 396 22499 424
rect 22527 396 22561 424
rect 22589 396 22623 424
rect 22651 396 22699 424
rect 22389 362 22699 396
rect 22389 334 22437 362
rect 22465 334 22499 362
rect 22527 334 22561 362
rect 22589 334 22623 362
rect 22651 334 22699 362
rect 22389 300 22699 334
rect 22389 272 22437 300
rect 22465 272 22499 300
rect 22527 272 22561 300
rect 22589 272 22623 300
rect 22651 272 22699 300
rect 22389 238 22699 272
rect 22389 210 22437 238
rect 22465 210 22499 238
rect 22527 210 22561 238
rect 22589 210 22623 238
rect 22651 210 22699 238
rect 22389 162 22699 210
rect 29529 20959 29839 29745
rect 29529 20931 29577 20959
rect 29605 20931 29639 20959
rect 29667 20931 29701 20959
rect 29729 20931 29763 20959
rect 29791 20931 29839 20959
rect 29529 20897 29839 20931
rect 29529 20869 29577 20897
rect 29605 20869 29639 20897
rect 29667 20869 29701 20897
rect 29729 20869 29763 20897
rect 29791 20869 29839 20897
rect 29529 20835 29839 20869
rect 29529 20807 29577 20835
rect 29605 20807 29639 20835
rect 29667 20807 29701 20835
rect 29729 20807 29763 20835
rect 29791 20807 29839 20835
rect 29529 20773 29839 20807
rect 29529 20745 29577 20773
rect 29605 20745 29639 20773
rect 29667 20745 29701 20773
rect 29729 20745 29763 20773
rect 29791 20745 29839 20773
rect 29529 11959 29839 20745
rect 29529 11931 29577 11959
rect 29605 11931 29639 11959
rect 29667 11931 29701 11959
rect 29729 11931 29763 11959
rect 29791 11931 29839 11959
rect 29529 11897 29839 11931
rect 29529 11869 29577 11897
rect 29605 11869 29639 11897
rect 29667 11869 29701 11897
rect 29729 11869 29763 11897
rect 29791 11869 29839 11897
rect 29529 11835 29839 11869
rect 29529 11807 29577 11835
rect 29605 11807 29639 11835
rect 29667 11807 29701 11835
rect 29729 11807 29763 11835
rect 29791 11807 29839 11835
rect 29529 11773 29839 11807
rect 29529 11745 29577 11773
rect 29605 11745 29639 11773
rect 29667 11745 29701 11773
rect 29729 11745 29763 11773
rect 29791 11745 29839 11773
rect 29529 2959 29839 11745
rect 29529 2931 29577 2959
rect 29605 2931 29639 2959
rect 29667 2931 29701 2959
rect 29729 2931 29763 2959
rect 29791 2931 29839 2959
rect 29529 2897 29839 2931
rect 29529 2869 29577 2897
rect 29605 2869 29639 2897
rect 29667 2869 29701 2897
rect 29729 2869 29763 2897
rect 29791 2869 29839 2897
rect 29529 2835 29839 2869
rect 29529 2807 29577 2835
rect 29605 2807 29639 2835
rect 29667 2807 29701 2835
rect 29729 2807 29763 2835
rect 29791 2807 29839 2835
rect 29529 2773 29839 2807
rect 29529 2745 29577 2773
rect 29605 2745 29639 2773
rect 29667 2745 29701 2773
rect 29729 2745 29763 2773
rect 29791 2745 29839 2773
rect 29529 904 29839 2745
rect 29529 876 29577 904
rect 29605 876 29639 904
rect 29667 876 29701 904
rect 29729 876 29763 904
rect 29791 876 29839 904
rect 29529 842 29839 876
rect 29529 814 29577 842
rect 29605 814 29639 842
rect 29667 814 29701 842
rect 29729 814 29763 842
rect 29791 814 29839 842
rect 29529 780 29839 814
rect 29529 752 29577 780
rect 29605 752 29639 780
rect 29667 752 29701 780
rect 29729 752 29763 780
rect 29791 752 29839 780
rect 29529 718 29839 752
rect 29529 690 29577 718
rect 29605 690 29639 718
rect 29667 690 29701 718
rect 29729 690 29763 718
rect 29791 690 29839 718
rect 29529 162 29839 690
rect 31389 299670 31699 299718
rect 31389 299642 31437 299670
rect 31465 299642 31499 299670
rect 31527 299642 31561 299670
rect 31589 299642 31623 299670
rect 31651 299642 31699 299670
rect 31389 299608 31699 299642
rect 31389 299580 31437 299608
rect 31465 299580 31499 299608
rect 31527 299580 31561 299608
rect 31589 299580 31623 299608
rect 31651 299580 31699 299608
rect 31389 299546 31699 299580
rect 31389 299518 31437 299546
rect 31465 299518 31499 299546
rect 31527 299518 31561 299546
rect 31589 299518 31623 299546
rect 31651 299518 31699 299546
rect 31389 299484 31699 299518
rect 31389 299456 31437 299484
rect 31465 299456 31499 299484
rect 31527 299456 31561 299484
rect 31589 299456 31623 299484
rect 31651 299456 31699 299484
rect 31389 293959 31699 299456
rect 31389 293931 31437 293959
rect 31465 293931 31499 293959
rect 31527 293931 31561 293959
rect 31589 293931 31623 293959
rect 31651 293931 31699 293959
rect 31389 293897 31699 293931
rect 31389 293869 31437 293897
rect 31465 293869 31499 293897
rect 31527 293869 31561 293897
rect 31589 293869 31623 293897
rect 31651 293869 31699 293897
rect 31389 293835 31699 293869
rect 31389 293807 31437 293835
rect 31465 293807 31499 293835
rect 31527 293807 31561 293835
rect 31589 293807 31623 293835
rect 31651 293807 31699 293835
rect 31389 293773 31699 293807
rect 31389 293745 31437 293773
rect 31465 293745 31499 293773
rect 31527 293745 31561 293773
rect 31589 293745 31623 293773
rect 31651 293745 31699 293773
rect 31389 284959 31699 293745
rect 31389 284931 31437 284959
rect 31465 284931 31499 284959
rect 31527 284931 31561 284959
rect 31589 284931 31623 284959
rect 31651 284931 31699 284959
rect 31389 284897 31699 284931
rect 31389 284869 31437 284897
rect 31465 284869 31499 284897
rect 31527 284869 31561 284897
rect 31589 284869 31623 284897
rect 31651 284869 31699 284897
rect 31389 284835 31699 284869
rect 31389 284807 31437 284835
rect 31465 284807 31499 284835
rect 31527 284807 31561 284835
rect 31589 284807 31623 284835
rect 31651 284807 31699 284835
rect 31389 284773 31699 284807
rect 31389 284745 31437 284773
rect 31465 284745 31499 284773
rect 31527 284745 31561 284773
rect 31589 284745 31623 284773
rect 31651 284745 31699 284773
rect 31389 275959 31699 284745
rect 31389 275931 31437 275959
rect 31465 275931 31499 275959
rect 31527 275931 31561 275959
rect 31589 275931 31623 275959
rect 31651 275931 31699 275959
rect 31389 275897 31699 275931
rect 31389 275869 31437 275897
rect 31465 275869 31499 275897
rect 31527 275869 31561 275897
rect 31589 275869 31623 275897
rect 31651 275869 31699 275897
rect 31389 275835 31699 275869
rect 31389 275807 31437 275835
rect 31465 275807 31499 275835
rect 31527 275807 31561 275835
rect 31589 275807 31623 275835
rect 31651 275807 31699 275835
rect 31389 275773 31699 275807
rect 31389 275745 31437 275773
rect 31465 275745 31499 275773
rect 31527 275745 31561 275773
rect 31589 275745 31623 275773
rect 31651 275745 31699 275773
rect 31389 266959 31699 275745
rect 31389 266931 31437 266959
rect 31465 266931 31499 266959
rect 31527 266931 31561 266959
rect 31589 266931 31623 266959
rect 31651 266931 31699 266959
rect 31389 266897 31699 266931
rect 31389 266869 31437 266897
rect 31465 266869 31499 266897
rect 31527 266869 31561 266897
rect 31589 266869 31623 266897
rect 31651 266869 31699 266897
rect 31389 266835 31699 266869
rect 31389 266807 31437 266835
rect 31465 266807 31499 266835
rect 31527 266807 31561 266835
rect 31589 266807 31623 266835
rect 31651 266807 31699 266835
rect 31389 266773 31699 266807
rect 31389 266745 31437 266773
rect 31465 266745 31499 266773
rect 31527 266745 31561 266773
rect 31589 266745 31623 266773
rect 31651 266745 31699 266773
rect 31389 257959 31699 266745
rect 31389 257931 31437 257959
rect 31465 257931 31499 257959
rect 31527 257931 31561 257959
rect 31589 257931 31623 257959
rect 31651 257931 31699 257959
rect 31389 257897 31699 257931
rect 31389 257869 31437 257897
rect 31465 257869 31499 257897
rect 31527 257869 31561 257897
rect 31589 257869 31623 257897
rect 31651 257869 31699 257897
rect 31389 257835 31699 257869
rect 31389 257807 31437 257835
rect 31465 257807 31499 257835
rect 31527 257807 31561 257835
rect 31589 257807 31623 257835
rect 31651 257807 31699 257835
rect 31389 257773 31699 257807
rect 31389 257745 31437 257773
rect 31465 257745 31499 257773
rect 31527 257745 31561 257773
rect 31589 257745 31623 257773
rect 31651 257745 31699 257773
rect 31389 248959 31699 257745
rect 38529 299190 38839 299718
rect 38529 299162 38577 299190
rect 38605 299162 38639 299190
rect 38667 299162 38701 299190
rect 38729 299162 38763 299190
rect 38791 299162 38839 299190
rect 38529 299128 38839 299162
rect 38529 299100 38577 299128
rect 38605 299100 38639 299128
rect 38667 299100 38701 299128
rect 38729 299100 38763 299128
rect 38791 299100 38839 299128
rect 38529 299066 38839 299100
rect 38529 299038 38577 299066
rect 38605 299038 38639 299066
rect 38667 299038 38701 299066
rect 38729 299038 38763 299066
rect 38791 299038 38839 299066
rect 38529 299004 38839 299038
rect 38529 298976 38577 299004
rect 38605 298976 38639 299004
rect 38667 298976 38701 299004
rect 38729 298976 38763 299004
rect 38791 298976 38839 299004
rect 38529 290959 38839 298976
rect 38529 290931 38577 290959
rect 38605 290931 38639 290959
rect 38667 290931 38701 290959
rect 38729 290931 38763 290959
rect 38791 290931 38839 290959
rect 38529 290897 38839 290931
rect 38529 290869 38577 290897
rect 38605 290869 38639 290897
rect 38667 290869 38701 290897
rect 38729 290869 38763 290897
rect 38791 290869 38839 290897
rect 38529 290835 38839 290869
rect 38529 290807 38577 290835
rect 38605 290807 38639 290835
rect 38667 290807 38701 290835
rect 38729 290807 38763 290835
rect 38791 290807 38839 290835
rect 38529 290773 38839 290807
rect 38529 290745 38577 290773
rect 38605 290745 38639 290773
rect 38667 290745 38701 290773
rect 38729 290745 38763 290773
rect 38791 290745 38839 290773
rect 38529 281959 38839 290745
rect 38529 281931 38577 281959
rect 38605 281931 38639 281959
rect 38667 281931 38701 281959
rect 38729 281931 38763 281959
rect 38791 281931 38839 281959
rect 38529 281897 38839 281931
rect 38529 281869 38577 281897
rect 38605 281869 38639 281897
rect 38667 281869 38701 281897
rect 38729 281869 38763 281897
rect 38791 281869 38839 281897
rect 38529 281835 38839 281869
rect 38529 281807 38577 281835
rect 38605 281807 38639 281835
rect 38667 281807 38701 281835
rect 38729 281807 38763 281835
rect 38791 281807 38839 281835
rect 38529 281773 38839 281807
rect 38529 281745 38577 281773
rect 38605 281745 38639 281773
rect 38667 281745 38701 281773
rect 38729 281745 38763 281773
rect 38791 281745 38839 281773
rect 38529 272959 38839 281745
rect 38529 272931 38577 272959
rect 38605 272931 38639 272959
rect 38667 272931 38701 272959
rect 38729 272931 38763 272959
rect 38791 272931 38839 272959
rect 38529 272897 38839 272931
rect 38529 272869 38577 272897
rect 38605 272869 38639 272897
rect 38667 272869 38701 272897
rect 38729 272869 38763 272897
rect 38791 272869 38839 272897
rect 38529 272835 38839 272869
rect 38529 272807 38577 272835
rect 38605 272807 38639 272835
rect 38667 272807 38701 272835
rect 38729 272807 38763 272835
rect 38791 272807 38839 272835
rect 38529 272773 38839 272807
rect 38529 272745 38577 272773
rect 38605 272745 38639 272773
rect 38667 272745 38701 272773
rect 38729 272745 38763 272773
rect 38791 272745 38839 272773
rect 38529 263959 38839 272745
rect 38529 263931 38577 263959
rect 38605 263931 38639 263959
rect 38667 263931 38701 263959
rect 38729 263931 38763 263959
rect 38791 263931 38839 263959
rect 38529 263897 38839 263931
rect 38529 263869 38577 263897
rect 38605 263869 38639 263897
rect 38667 263869 38701 263897
rect 38729 263869 38763 263897
rect 38791 263869 38839 263897
rect 38529 263835 38839 263869
rect 38529 263807 38577 263835
rect 38605 263807 38639 263835
rect 38667 263807 38701 263835
rect 38729 263807 38763 263835
rect 38791 263807 38839 263835
rect 38529 263773 38839 263807
rect 38529 263745 38577 263773
rect 38605 263745 38639 263773
rect 38667 263745 38701 263773
rect 38729 263745 38763 263773
rect 38791 263745 38839 263773
rect 38529 254959 38839 263745
rect 38529 254931 38577 254959
rect 38605 254931 38639 254959
rect 38667 254931 38701 254959
rect 38729 254931 38763 254959
rect 38791 254931 38839 254959
rect 38529 254897 38839 254931
rect 38529 254869 38577 254897
rect 38605 254869 38639 254897
rect 38667 254869 38701 254897
rect 38729 254869 38763 254897
rect 38791 254869 38839 254897
rect 38529 254835 38839 254869
rect 38529 254807 38577 254835
rect 38605 254807 38639 254835
rect 38667 254807 38701 254835
rect 38729 254807 38763 254835
rect 38791 254807 38839 254835
rect 38529 254773 38839 254807
rect 38529 254745 38577 254773
rect 38605 254745 38639 254773
rect 38667 254745 38701 254773
rect 38729 254745 38763 254773
rect 38791 254745 38839 254773
rect 38529 254075 38839 254745
rect 40389 299670 40699 299718
rect 40389 299642 40437 299670
rect 40465 299642 40499 299670
rect 40527 299642 40561 299670
rect 40589 299642 40623 299670
rect 40651 299642 40699 299670
rect 40389 299608 40699 299642
rect 40389 299580 40437 299608
rect 40465 299580 40499 299608
rect 40527 299580 40561 299608
rect 40589 299580 40623 299608
rect 40651 299580 40699 299608
rect 40389 299546 40699 299580
rect 40389 299518 40437 299546
rect 40465 299518 40499 299546
rect 40527 299518 40561 299546
rect 40589 299518 40623 299546
rect 40651 299518 40699 299546
rect 40389 299484 40699 299518
rect 40389 299456 40437 299484
rect 40465 299456 40499 299484
rect 40527 299456 40561 299484
rect 40589 299456 40623 299484
rect 40651 299456 40699 299484
rect 40389 293959 40699 299456
rect 40389 293931 40437 293959
rect 40465 293931 40499 293959
rect 40527 293931 40561 293959
rect 40589 293931 40623 293959
rect 40651 293931 40699 293959
rect 40389 293897 40699 293931
rect 40389 293869 40437 293897
rect 40465 293869 40499 293897
rect 40527 293869 40561 293897
rect 40589 293869 40623 293897
rect 40651 293869 40699 293897
rect 40389 293835 40699 293869
rect 40389 293807 40437 293835
rect 40465 293807 40499 293835
rect 40527 293807 40561 293835
rect 40589 293807 40623 293835
rect 40651 293807 40699 293835
rect 40389 293773 40699 293807
rect 40389 293745 40437 293773
rect 40465 293745 40499 293773
rect 40527 293745 40561 293773
rect 40589 293745 40623 293773
rect 40651 293745 40699 293773
rect 40389 284959 40699 293745
rect 40389 284931 40437 284959
rect 40465 284931 40499 284959
rect 40527 284931 40561 284959
rect 40589 284931 40623 284959
rect 40651 284931 40699 284959
rect 40389 284897 40699 284931
rect 40389 284869 40437 284897
rect 40465 284869 40499 284897
rect 40527 284869 40561 284897
rect 40589 284869 40623 284897
rect 40651 284869 40699 284897
rect 40389 284835 40699 284869
rect 40389 284807 40437 284835
rect 40465 284807 40499 284835
rect 40527 284807 40561 284835
rect 40589 284807 40623 284835
rect 40651 284807 40699 284835
rect 40389 284773 40699 284807
rect 40389 284745 40437 284773
rect 40465 284745 40499 284773
rect 40527 284745 40561 284773
rect 40589 284745 40623 284773
rect 40651 284745 40699 284773
rect 40389 275959 40699 284745
rect 40389 275931 40437 275959
rect 40465 275931 40499 275959
rect 40527 275931 40561 275959
rect 40589 275931 40623 275959
rect 40651 275931 40699 275959
rect 40389 275897 40699 275931
rect 40389 275869 40437 275897
rect 40465 275869 40499 275897
rect 40527 275869 40561 275897
rect 40589 275869 40623 275897
rect 40651 275869 40699 275897
rect 40389 275835 40699 275869
rect 40389 275807 40437 275835
rect 40465 275807 40499 275835
rect 40527 275807 40561 275835
rect 40589 275807 40623 275835
rect 40651 275807 40699 275835
rect 40389 275773 40699 275807
rect 40389 275745 40437 275773
rect 40465 275745 40499 275773
rect 40527 275745 40561 275773
rect 40589 275745 40623 275773
rect 40651 275745 40699 275773
rect 40389 266959 40699 275745
rect 40389 266931 40437 266959
rect 40465 266931 40499 266959
rect 40527 266931 40561 266959
rect 40589 266931 40623 266959
rect 40651 266931 40699 266959
rect 40389 266897 40699 266931
rect 40389 266869 40437 266897
rect 40465 266869 40499 266897
rect 40527 266869 40561 266897
rect 40589 266869 40623 266897
rect 40651 266869 40699 266897
rect 40389 266835 40699 266869
rect 40389 266807 40437 266835
rect 40465 266807 40499 266835
rect 40527 266807 40561 266835
rect 40589 266807 40623 266835
rect 40651 266807 40699 266835
rect 40389 266773 40699 266807
rect 40389 266745 40437 266773
rect 40465 266745 40499 266773
rect 40527 266745 40561 266773
rect 40589 266745 40623 266773
rect 40651 266745 40699 266773
rect 40389 257959 40699 266745
rect 40389 257931 40437 257959
rect 40465 257931 40499 257959
rect 40527 257931 40561 257959
rect 40589 257931 40623 257959
rect 40651 257931 40699 257959
rect 40389 257897 40699 257931
rect 40389 257869 40437 257897
rect 40465 257869 40499 257897
rect 40527 257869 40561 257897
rect 40589 257869 40623 257897
rect 40651 257869 40699 257897
rect 40389 257835 40699 257869
rect 40389 257807 40437 257835
rect 40465 257807 40499 257835
rect 40527 257807 40561 257835
rect 40589 257807 40623 257835
rect 40651 257807 40699 257835
rect 40389 257773 40699 257807
rect 40389 257745 40437 257773
rect 40465 257745 40499 257773
rect 40527 257745 40561 257773
rect 40589 257745 40623 257773
rect 40651 257745 40699 257773
rect 40389 254394 40699 257745
rect 47529 299190 47839 299718
rect 47529 299162 47577 299190
rect 47605 299162 47639 299190
rect 47667 299162 47701 299190
rect 47729 299162 47763 299190
rect 47791 299162 47839 299190
rect 47529 299128 47839 299162
rect 47529 299100 47577 299128
rect 47605 299100 47639 299128
rect 47667 299100 47701 299128
rect 47729 299100 47763 299128
rect 47791 299100 47839 299128
rect 47529 299066 47839 299100
rect 47529 299038 47577 299066
rect 47605 299038 47639 299066
rect 47667 299038 47701 299066
rect 47729 299038 47763 299066
rect 47791 299038 47839 299066
rect 47529 299004 47839 299038
rect 47529 298976 47577 299004
rect 47605 298976 47639 299004
rect 47667 298976 47701 299004
rect 47729 298976 47763 299004
rect 47791 298976 47839 299004
rect 47529 290959 47839 298976
rect 47529 290931 47577 290959
rect 47605 290931 47639 290959
rect 47667 290931 47701 290959
rect 47729 290931 47763 290959
rect 47791 290931 47839 290959
rect 47529 290897 47839 290931
rect 47529 290869 47577 290897
rect 47605 290869 47639 290897
rect 47667 290869 47701 290897
rect 47729 290869 47763 290897
rect 47791 290869 47839 290897
rect 47529 290835 47839 290869
rect 47529 290807 47577 290835
rect 47605 290807 47639 290835
rect 47667 290807 47701 290835
rect 47729 290807 47763 290835
rect 47791 290807 47839 290835
rect 47529 290773 47839 290807
rect 47529 290745 47577 290773
rect 47605 290745 47639 290773
rect 47667 290745 47701 290773
rect 47729 290745 47763 290773
rect 47791 290745 47839 290773
rect 47529 281959 47839 290745
rect 47529 281931 47577 281959
rect 47605 281931 47639 281959
rect 47667 281931 47701 281959
rect 47729 281931 47763 281959
rect 47791 281931 47839 281959
rect 47529 281897 47839 281931
rect 47529 281869 47577 281897
rect 47605 281869 47639 281897
rect 47667 281869 47701 281897
rect 47729 281869 47763 281897
rect 47791 281869 47839 281897
rect 47529 281835 47839 281869
rect 47529 281807 47577 281835
rect 47605 281807 47639 281835
rect 47667 281807 47701 281835
rect 47729 281807 47763 281835
rect 47791 281807 47839 281835
rect 47529 281773 47839 281807
rect 47529 281745 47577 281773
rect 47605 281745 47639 281773
rect 47667 281745 47701 281773
rect 47729 281745 47763 281773
rect 47791 281745 47839 281773
rect 47529 272959 47839 281745
rect 47529 272931 47577 272959
rect 47605 272931 47639 272959
rect 47667 272931 47701 272959
rect 47729 272931 47763 272959
rect 47791 272931 47839 272959
rect 47529 272897 47839 272931
rect 47529 272869 47577 272897
rect 47605 272869 47639 272897
rect 47667 272869 47701 272897
rect 47729 272869 47763 272897
rect 47791 272869 47839 272897
rect 47529 272835 47839 272869
rect 47529 272807 47577 272835
rect 47605 272807 47639 272835
rect 47667 272807 47701 272835
rect 47729 272807 47763 272835
rect 47791 272807 47839 272835
rect 47529 272773 47839 272807
rect 47529 272745 47577 272773
rect 47605 272745 47639 272773
rect 47667 272745 47701 272773
rect 47729 272745 47763 272773
rect 47791 272745 47839 272773
rect 47529 263959 47839 272745
rect 47529 263931 47577 263959
rect 47605 263931 47639 263959
rect 47667 263931 47701 263959
rect 47729 263931 47763 263959
rect 47791 263931 47839 263959
rect 47529 263897 47839 263931
rect 47529 263869 47577 263897
rect 47605 263869 47639 263897
rect 47667 263869 47701 263897
rect 47729 263869 47763 263897
rect 47791 263869 47839 263897
rect 47529 263835 47839 263869
rect 47529 263807 47577 263835
rect 47605 263807 47639 263835
rect 47667 263807 47701 263835
rect 47729 263807 47763 263835
rect 47791 263807 47839 263835
rect 47529 263773 47839 263807
rect 47529 263745 47577 263773
rect 47605 263745 47639 263773
rect 47667 263745 47701 263773
rect 47729 263745 47763 263773
rect 47791 263745 47839 263773
rect 47529 254959 47839 263745
rect 47529 254931 47577 254959
rect 47605 254931 47639 254959
rect 47667 254931 47701 254959
rect 47729 254931 47763 254959
rect 47791 254931 47839 254959
rect 47529 254897 47839 254931
rect 47529 254869 47577 254897
rect 47605 254869 47639 254897
rect 47667 254869 47701 254897
rect 47729 254869 47763 254897
rect 47791 254869 47839 254897
rect 47529 254835 47839 254869
rect 47529 254807 47577 254835
rect 47605 254807 47639 254835
rect 47667 254807 47701 254835
rect 47729 254807 47763 254835
rect 47791 254807 47839 254835
rect 47529 254773 47839 254807
rect 47529 254745 47577 254773
rect 47605 254745 47639 254773
rect 47667 254745 47701 254773
rect 47729 254745 47763 254773
rect 47791 254745 47839 254773
rect 47529 254075 47839 254745
rect 49389 299670 49699 299718
rect 49389 299642 49437 299670
rect 49465 299642 49499 299670
rect 49527 299642 49561 299670
rect 49589 299642 49623 299670
rect 49651 299642 49699 299670
rect 49389 299608 49699 299642
rect 49389 299580 49437 299608
rect 49465 299580 49499 299608
rect 49527 299580 49561 299608
rect 49589 299580 49623 299608
rect 49651 299580 49699 299608
rect 49389 299546 49699 299580
rect 49389 299518 49437 299546
rect 49465 299518 49499 299546
rect 49527 299518 49561 299546
rect 49589 299518 49623 299546
rect 49651 299518 49699 299546
rect 49389 299484 49699 299518
rect 49389 299456 49437 299484
rect 49465 299456 49499 299484
rect 49527 299456 49561 299484
rect 49589 299456 49623 299484
rect 49651 299456 49699 299484
rect 49389 293959 49699 299456
rect 49389 293931 49437 293959
rect 49465 293931 49499 293959
rect 49527 293931 49561 293959
rect 49589 293931 49623 293959
rect 49651 293931 49699 293959
rect 49389 293897 49699 293931
rect 49389 293869 49437 293897
rect 49465 293869 49499 293897
rect 49527 293869 49561 293897
rect 49589 293869 49623 293897
rect 49651 293869 49699 293897
rect 49389 293835 49699 293869
rect 49389 293807 49437 293835
rect 49465 293807 49499 293835
rect 49527 293807 49561 293835
rect 49589 293807 49623 293835
rect 49651 293807 49699 293835
rect 49389 293773 49699 293807
rect 49389 293745 49437 293773
rect 49465 293745 49499 293773
rect 49527 293745 49561 293773
rect 49589 293745 49623 293773
rect 49651 293745 49699 293773
rect 49389 284959 49699 293745
rect 49389 284931 49437 284959
rect 49465 284931 49499 284959
rect 49527 284931 49561 284959
rect 49589 284931 49623 284959
rect 49651 284931 49699 284959
rect 49389 284897 49699 284931
rect 49389 284869 49437 284897
rect 49465 284869 49499 284897
rect 49527 284869 49561 284897
rect 49589 284869 49623 284897
rect 49651 284869 49699 284897
rect 49389 284835 49699 284869
rect 49389 284807 49437 284835
rect 49465 284807 49499 284835
rect 49527 284807 49561 284835
rect 49589 284807 49623 284835
rect 49651 284807 49699 284835
rect 49389 284773 49699 284807
rect 49389 284745 49437 284773
rect 49465 284745 49499 284773
rect 49527 284745 49561 284773
rect 49589 284745 49623 284773
rect 49651 284745 49699 284773
rect 49389 275959 49699 284745
rect 49389 275931 49437 275959
rect 49465 275931 49499 275959
rect 49527 275931 49561 275959
rect 49589 275931 49623 275959
rect 49651 275931 49699 275959
rect 49389 275897 49699 275931
rect 49389 275869 49437 275897
rect 49465 275869 49499 275897
rect 49527 275869 49561 275897
rect 49589 275869 49623 275897
rect 49651 275869 49699 275897
rect 49389 275835 49699 275869
rect 49389 275807 49437 275835
rect 49465 275807 49499 275835
rect 49527 275807 49561 275835
rect 49589 275807 49623 275835
rect 49651 275807 49699 275835
rect 49389 275773 49699 275807
rect 49389 275745 49437 275773
rect 49465 275745 49499 275773
rect 49527 275745 49561 275773
rect 49589 275745 49623 275773
rect 49651 275745 49699 275773
rect 49389 266959 49699 275745
rect 49389 266931 49437 266959
rect 49465 266931 49499 266959
rect 49527 266931 49561 266959
rect 49589 266931 49623 266959
rect 49651 266931 49699 266959
rect 49389 266897 49699 266931
rect 49389 266869 49437 266897
rect 49465 266869 49499 266897
rect 49527 266869 49561 266897
rect 49589 266869 49623 266897
rect 49651 266869 49699 266897
rect 49389 266835 49699 266869
rect 49389 266807 49437 266835
rect 49465 266807 49499 266835
rect 49527 266807 49561 266835
rect 49589 266807 49623 266835
rect 49651 266807 49699 266835
rect 49389 266773 49699 266807
rect 49389 266745 49437 266773
rect 49465 266745 49499 266773
rect 49527 266745 49561 266773
rect 49589 266745 49623 266773
rect 49651 266745 49699 266773
rect 49389 257959 49699 266745
rect 49389 257931 49437 257959
rect 49465 257931 49499 257959
rect 49527 257931 49561 257959
rect 49589 257931 49623 257959
rect 49651 257931 49699 257959
rect 49389 257897 49699 257931
rect 49389 257869 49437 257897
rect 49465 257869 49499 257897
rect 49527 257869 49561 257897
rect 49589 257869 49623 257897
rect 49651 257869 49699 257897
rect 49389 257835 49699 257869
rect 49389 257807 49437 257835
rect 49465 257807 49499 257835
rect 49527 257807 49561 257835
rect 49589 257807 49623 257835
rect 49651 257807 49699 257835
rect 49389 257773 49699 257807
rect 49389 257745 49437 257773
rect 49465 257745 49499 257773
rect 49527 257745 49561 257773
rect 49589 257745 49623 257773
rect 49651 257745 49699 257773
rect 49389 254075 49699 257745
rect 56529 299190 56839 299718
rect 56529 299162 56577 299190
rect 56605 299162 56639 299190
rect 56667 299162 56701 299190
rect 56729 299162 56763 299190
rect 56791 299162 56839 299190
rect 56529 299128 56839 299162
rect 56529 299100 56577 299128
rect 56605 299100 56639 299128
rect 56667 299100 56701 299128
rect 56729 299100 56763 299128
rect 56791 299100 56839 299128
rect 56529 299066 56839 299100
rect 56529 299038 56577 299066
rect 56605 299038 56639 299066
rect 56667 299038 56701 299066
rect 56729 299038 56763 299066
rect 56791 299038 56839 299066
rect 56529 299004 56839 299038
rect 56529 298976 56577 299004
rect 56605 298976 56639 299004
rect 56667 298976 56701 299004
rect 56729 298976 56763 299004
rect 56791 298976 56839 299004
rect 56529 290959 56839 298976
rect 56529 290931 56577 290959
rect 56605 290931 56639 290959
rect 56667 290931 56701 290959
rect 56729 290931 56763 290959
rect 56791 290931 56839 290959
rect 56529 290897 56839 290931
rect 56529 290869 56577 290897
rect 56605 290869 56639 290897
rect 56667 290869 56701 290897
rect 56729 290869 56763 290897
rect 56791 290869 56839 290897
rect 56529 290835 56839 290869
rect 56529 290807 56577 290835
rect 56605 290807 56639 290835
rect 56667 290807 56701 290835
rect 56729 290807 56763 290835
rect 56791 290807 56839 290835
rect 56529 290773 56839 290807
rect 56529 290745 56577 290773
rect 56605 290745 56639 290773
rect 56667 290745 56701 290773
rect 56729 290745 56763 290773
rect 56791 290745 56839 290773
rect 56529 281959 56839 290745
rect 56529 281931 56577 281959
rect 56605 281931 56639 281959
rect 56667 281931 56701 281959
rect 56729 281931 56763 281959
rect 56791 281931 56839 281959
rect 56529 281897 56839 281931
rect 56529 281869 56577 281897
rect 56605 281869 56639 281897
rect 56667 281869 56701 281897
rect 56729 281869 56763 281897
rect 56791 281869 56839 281897
rect 56529 281835 56839 281869
rect 56529 281807 56577 281835
rect 56605 281807 56639 281835
rect 56667 281807 56701 281835
rect 56729 281807 56763 281835
rect 56791 281807 56839 281835
rect 56529 281773 56839 281807
rect 56529 281745 56577 281773
rect 56605 281745 56639 281773
rect 56667 281745 56701 281773
rect 56729 281745 56763 281773
rect 56791 281745 56839 281773
rect 56529 272959 56839 281745
rect 56529 272931 56577 272959
rect 56605 272931 56639 272959
rect 56667 272931 56701 272959
rect 56729 272931 56763 272959
rect 56791 272931 56839 272959
rect 56529 272897 56839 272931
rect 56529 272869 56577 272897
rect 56605 272869 56639 272897
rect 56667 272869 56701 272897
rect 56729 272869 56763 272897
rect 56791 272869 56839 272897
rect 56529 272835 56839 272869
rect 56529 272807 56577 272835
rect 56605 272807 56639 272835
rect 56667 272807 56701 272835
rect 56729 272807 56763 272835
rect 56791 272807 56839 272835
rect 56529 272773 56839 272807
rect 56529 272745 56577 272773
rect 56605 272745 56639 272773
rect 56667 272745 56701 272773
rect 56729 272745 56763 272773
rect 56791 272745 56839 272773
rect 56529 263959 56839 272745
rect 56529 263931 56577 263959
rect 56605 263931 56639 263959
rect 56667 263931 56701 263959
rect 56729 263931 56763 263959
rect 56791 263931 56839 263959
rect 56529 263897 56839 263931
rect 56529 263869 56577 263897
rect 56605 263869 56639 263897
rect 56667 263869 56701 263897
rect 56729 263869 56763 263897
rect 56791 263869 56839 263897
rect 56529 263835 56839 263869
rect 56529 263807 56577 263835
rect 56605 263807 56639 263835
rect 56667 263807 56701 263835
rect 56729 263807 56763 263835
rect 56791 263807 56839 263835
rect 56529 263773 56839 263807
rect 56529 263745 56577 263773
rect 56605 263745 56639 263773
rect 56667 263745 56701 263773
rect 56729 263745 56763 263773
rect 56791 263745 56839 263773
rect 56529 254959 56839 263745
rect 56529 254931 56577 254959
rect 56605 254931 56639 254959
rect 56667 254931 56701 254959
rect 56729 254931 56763 254959
rect 56791 254931 56839 254959
rect 56529 254897 56839 254931
rect 56529 254869 56577 254897
rect 56605 254869 56639 254897
rect 56667 254869 56701 254897
rect 56729 254869 56763 254897
rect 56791 254869 56839 254897
rect 56529 254835 56839 254869
rect 56529 254807 56577 254835
rect 56605 254807 56639 254835
rect 56667 254807 56701 254835
rect 56729 254807 56763 254835
rect 56791 254807 56839 254835
rect 56529 254773 56839 254807
rect 56529 254745 56577 254773
rect 56605 254745 56639 254773
rect 56667 254745 56701 254773
rect 56729 254745 56763 254773
rect 56791 254745 56839 254773
rect 56529 254075 56839 254745
rect 58389 299670 58699 299718
rect 58389 299642 58437 299670
rect 58465 299642 58499 299670
rect 58527 299642 58561 299670
rect 58589 299642 58623 299670
rect 58651 299642 58699 299670
rect 58389 299608 58699 299642
rect 58389 299580 58437 299608
rect 58465 299580 58499 299608
rect 58527 299580 58561 299608
rect 58589 299580 58623 299608
rect 58651 299580 58699 299608
rect 58389 299546 58699 299580
rect 58389 299518 58437 299546
rect 58465 299518 58499 299546
rect 58527 299518 58561 299546
rect 58589 299518 58623 299546
rect 58651 299518 58699 299546
rect 58389 299484 58699 299518
rect 58389 299456 58437 299484
rect 58465 299456 58499 299484
rect 58527 299456 58561 299484
rect 58589 299456 58623 299484
rect 58651 299456 58699 299484
rect 58389 293959 58699 299456
rect 58389 293931 58437 293959
rect 58465 293931 58499 293959
rect 58527 293931 58561 293959
rect 58589 293931 58623 293959
rect 58651 293931 58699 293959
rect 58389 293897 58699 293931
rect 58389 293869 58437 293897
rect 58465 293869 58499 293897
rect 58527 293869 58561 293897
rect 58589 293869 58623 293897
rect 58651 293869 58699 293897
rect 58389 293835 58699 293869
rect 58389 293807 58437 293835
rect 58465 293807 58499 293835
rect 58527 293807 58561 293835
rect 58589 293807 58623 293835
rect 58651 293807 58699 293835
rect 58389 293773 58699 293807
rect 58389 293745 58437 293773
rect 58465 293745 58499 293773
rect 58527 293745 58561 293773
rect 58589 293745 58623 293773
rect 58651 293745 58699 293773
rect 58389 284959 58699 293745
rect 58389 284931 58437 284959
rect 58465 284931 58499 284959
rect 58527 284931 58561 284959
rect 58589 284931 58623 284959
rect 58651 284931 58699 284959
rect 58389 284897 58699 284931
rect 58389 284869 58437 284897
rect 58465 284869 58499 284897
rect 58527 284869 58561 284897
rect 58589 284869 58623 284897
rect 58651 284869 58699 284897
rect 58389 284835 58699 284869
rect 58389 284807 58437 284835
rect 58465 284807 58499 284835
rect 58527 284807 58561 284835
rect 58589 284807 58623 284835
rect 58651 284807 58699 284835
rect 58389 284773 58699 284807
rect 58389 284745 58437 284773
rect 58465 284745 58499 284773
rect 58527 284745 58561 284773
rect 58589 284745 58623 284773
rect 58651 284745 58699 284773
rect 58389 275959 58699 284745
rect 58389 275931 58437 275959
rect 58465 275931 58499 275959
rect 58527 275931 58561 275959
rect 58589 275931 58623 275959
rect 58651 275931 58699 275959
rect 58389 275897 58699 275931
rect 58389 275869 58437 275897
rect 58465 275869 58499 275897
rect 58527 275869 58561 275897
rect 58589 275869 58623 275897
rect 58651 275869 58699 275897
rect 58389 275835 58699 275869
rect 58389 275807 58437 275835
rect 58465 275807 58499 275835
rect 58527 275807 58561 275835
rect 58589 275807 58623 275835
rect 58651 275807 58699 275835
rect 58389 275773 58699 275807
rect 58389 275745 58437 275773
rect 58465 275745 58499 275773
rect 58527 275745 58561 275773
rect 58589 275745 58623 275773
rect 58651 275745 58699 275773
rect 58389 266959 58699 275745
rect 58389 266931 58437 266959
rect 58465 266931 58499 266959
rect 58527 266931 58561 266959
rect 58589 266931 58623 266959
rect 58651 266931 58699 266959
rect 58389 266897 58699 266931
rect 58389 266869 58437 266897
rect 58465 266869 58499 266897
rect 58527 266869 58561 266897
rect 58589 266869 58623 266897
rect 58651 266869 58699 266897
rect 58389 266835 58699 266869
rect 58389 266807 58437 266835
rect 58465 266807 58499 266835
rect 58527 266807 58561 266835
rect 58589 266807 58623 266835
rect 58651 266807 58699 266835
rect 58389 266773 58699 266807
rect 58389 266745 58437 266773
rect 58465 266745 58499 266773
rect 58527 266745 58561 266773
rect 58589 266745 58623 266773
rect 58651 266745 58699 266773
rect 58389 257959 58699 266745
rect 58389 257931 58437 257959
rect 58465 257931 58499 257959
rect 58527 257931 58561 257959
rect 58589 257931 58623 257959
rect 58651 257931 58699 257959
rect 58389 257897 58699 257931
rect 58389 257869 58437 257897
rect 58465 257869 58499 257897
rect 58527 257869 58561 257897
rect 58589 257869 58623 257897
rect 58651 257869 58699 257897
rect 58389 257835 58699 257869
rect 58389 257807 58437 257835
rect 58465 257807 58499 257835
rect 58527 257807 58561 257835
rect 58589 257807 58623 257835
rect 58651 257807 58699 257835
rect 58389 257773 58699 257807
rect 58389 257745 58437 257773
rect 58465 257745 58499 257773
rect 58527 257745 58561 257773
rect 58589 257745 58623 257773
rect 58651 257745 58699 257773
rect 58389 254075 58699 257745
rect 65529 299190 65839 299718
rect 65529 299162 65577 299190
rect 65605 299162 65639 299190
rect 65667 299162 65701 299190
rect 65729 299162 65763 299190
rect 65791 299162 65839 299190
rect 65529 299128 65839 299162
rect 65529 299100 65577 299128
rect 65605 299100 65639 299128
rect 65667 299100 65701 299128
rect 65729 299100 65763 299128
rect 65791 299100 65839 299128
rect 65529 299066 65839 299100
rect 65529 299038 65577 299066
rect 65605 299038 65639 299066
rect 65667 299038 65701 299066
rect 65729 299038 65763 299066
rect 65791 299038 65839 299066
rect 65529 299004 65839 299038
rect 65529 298976 65577 299004
rect 65605 298976 65639 299004
rect 65667 298976 65701 299004
rect 65729 298976 65763 299004
rect 65791 298976 65839 299004
rect 65529 290959 65839 298976
rect 65529 290931 65577 290959
rect 65605 290931 65639 290959
rect 65667 290931 65701 290959
rect 65729 290931 65763 290959
rect 65791 290931 65839 290959
rect 65529 290897 65839 290931
rect 65529 290869 65577 290897
rect 65605 290869 65639 290897
rect 65667 290869 65701 290897
rect 65729 290869 65763 290897
rect 65791 290869 65839 290897
rect 65529 290835 65839 290869
rect 65529 290807 65577 290835
rect 65605 290807 65639 290835
rect 65667 290807 65701 290835
rect 65729 290807 65763 290835
rect 65791 290807 65839 290835
rect 65529 290773 65839 290807
rect 65529 290745 65577 290773
rect 65605 290745 65639 290773
rect 65667 290745 65701 290773
rect 65729 290745 65763 290773
rect 65791 290745 65839 290773
rect 65529 281959 65839 290745
rect 65529 281931 65577 281959
rect 65605 281931 65639 281959
rect 65667 281931 65701 281959
rect 65729 281931 65763 281959
rect 65791 281931 65839 281959
rect 65529 281897 65839 281931
rect 65529 281869 65577 281897
rect 65605 281869 65639 281897
rect 65667 281869 65701 281897
rect 65729 281869 65763 281897
rect 65791 281869 65839 281897
rect 65529 281835 65839 281869
rect 65529 281807 65577 281835
rect 65605 281807 65639 281835
rect 65667 281807 65701 281835
rect 65729 281807 65763 281835
rect 65791 281807 65839 281835
rect 65529 281773 65839 281807
rect 65529 281745 65577 281773
rect 65605 281745 65639 281773
rect 65667 281745 65701 281773
rect 65729 281745 65763 281773
rect 65791 281745 65839 281773
rect 65529 272959 65839 281745
rect 65529 272931 65577 272959
rect 65605 272931 65639 272959
rect 65667 272931 65701 272959
rect 65729 272931 65763 272959
rect 65791 272931 65839 272959
rect 65529 272897 65839 272931
rect 65529 272869 65577 272897
rect 65605 272869 65639 272897
rect 65667 272869 65701 272897
rect 65729 272869 65763 272897
rect 65791 272869 65839 272897
rect 65529 272835 65839 272869
rect 65529 272807 65577 272835
rect 65605 272807 65639 272835
rect 65667 272807 65701 272835
rect 65729 272807 65763 272835
rect 65791 272807 65839 272835
rect 65529 272773 65839 272807
rect 65529 272745 65577 272773
rect 65605 272745 65639 272773
rect 65667 272745 65701 272773
rect 65729 272745 65763 272773
rect 65791 272745 65839 272773
rect 65529 263959 65839 272745
rect 65529 263931 65577 263959
rect 65605 263931 65639 263959
rect 65667 263931 65701 263959
rect 65729 263931 65763 263959
rect 65791 263931 65839 263959
rect 65529 263897 65839 263931
rect 65529 263869 65577 263897
rect 65605 263869 65639 263897
rect 65667 263869 65701 263897
rect 65729 263869 65763 263897
rect 65791 263869 65839 263897
rect 65529 263835 65839 263869
rect 65529 263807 65577 263835
rect 65605 263807 65639 263835
rect 65667 263807 65701 263835
rect 65729 263807 65763 263835
rect 65791 263807 65839 263835
rect 65529 263773 65839 263807
rect 65529 263745 65577 263773
rect 65605 263745 65639 263773
rect 65667 263745 65701 263773
rect 65729 263745 65763 263773
rect 65791 263745 65839 263773
rect 65529 254959 65839 263745
rect 65529 254931 65577 254959
rect 65605 254931 65639 254959
rect 65667 254931 65701 254959
rect 65729 254931 65763 254959
rect 65791 254931 65839 254959
rect 65529 254897 65839 254931
rect 65529 254869 65577 254897
rect 65605 254869 65639 254897
rect 65667 254869 65701 254897
rect 65729 254869 65763 254897
rect 65791 254869 65839 254897
rect 65529 254835 65839 254869
rect 65529 254807 65577 254835
rect 65605 254807 65639 254835
rect 65667 254807 65701 254835
rect 65729 254807 65763 254835
rect 65791 254807 65839 254835
rect 65529 254773 65839 254807
rect 65529 254745 65577 254773
rect 65605 254745 65639 254773
rect 65667 254745 65701 254773
rect 65729 254745 65763 254773
rect 65791 254745 65839 254773
rect 65529 254075 65839 254745
rect 67389 299670 67699 299718
rect 67389 299642 67437 299670
rect 67465 299642 67499 299670
rect 67527 299642 67561 299670
rect 67589 299642 67623 299670
rect 67651 299642 67699 299670
rect 67389 299608 67699 299642
rect 67389 299580 67437 299608
rect 67465 299580 67499 299608
rect 67527 299580 67561 299608
rect 67589 299580 67623 299608
rect 67651 299580 67699 299608
rect 67389 299546 67699 299580
rect 67389 299518 67437 299546
rect 67465 299518 67499 299546
rect 67527 299518 67561 299546
rect 67589 299518 67623 299546
rect 67651 299518 67699 299546
rect 67389 299484 67699 299518
rect 67389 299456 67437 299484
rect 67465 299456 67499 299484
rect 67527 299456 67561 299484
rect 67589 299456 67623 299484
rect 67651 299456 67699 299484
rect 67389 293959 67699 299456
rect 67389 293931 67437 293959
rect 67465 293931 67499 293959
rect 67527 293931 67561 293959
rect 67589 293931 67623 293959
rect 67651 293931 67699 293959
rect 67389 293897 67699 293931
rect 67389 293869 67437 293897
rect 67465 293869 67499 293897
rect 67527 293869 67561 293897
rect 67589 293869 67623 293897
rect 67651 293869 67699 293897
rect 67389 293835 67699 293869
rect 67389 293807 67437 293835
rect 67465 293807 67499 293835
rect 67527 293807 67561 293835
rect 67589 293807 67623 293835
rect 67651 293807 67699 293835
rect 67389 293773 67699 293807
rect 67389 293745 67437 293773
rect 67465 293745 67499 293773
rect 67527 293745 67561 293773
rect 67589 293745 67623 293773
rect 67651 293745 67699 293773
rect 67389 284959 67699 293745
rect 67389 284931 67437 284959
rect 67465 284931 67499 284959
rect 67527 284931 67561 284959
rect 67589 284931 67623 284959
rect 67651 284931 67699 284959
rect 67389 284897 67699 284931
rect 67389 284869 67437 284897
rect 67465 284869 67499 284897
rect 67527 284869 67561 284897
rect 67589 284869 67623 284897
rect 67651 284869 67699 284897
rect 67389 284835 67699 284869
rect 67389 284807 67437 284835
rect 67465 284807 67499 284835
rect 67527 284807 67561 284835
rect 67589 284807 67623 284835
rect 67651 284807 67699 284835
rect 67389 284773 67699 284807
rect 67389 284745 67437 284773
rect 67465 284745 67499 284773
rect 67527 284745 67561 284773
rect 67589 284745 67623 284773
rect 67651 284745 67699 284773
rect 67389 275959 67699 284745
rect 67389 275931 67437 275959
rect 67465 275931 67499 275959
rect 67527 275931 67561 275959
rect 67589 275931 67623 275959
rect 67651 275931 67699 275959
rect 67389 275897 67699 275931
rect 67389 275869 67437 275897
rect 67465 275869 67499 275897
rect 67527 275869 67561 275897
rect 67589 275869 67623 275897
rect 67651 275869 67699 275897
rect 67389 275835 67699 275869
rect 67389 275807 67437 275835
rect 67465 275807 67499 275835
rect 67527 275807 67561 275835
rect 67589 275807 67623 275835
rect 67651 275807 67699 275835
rect 67389 275773 67699 275807
rect 67389 275745 67437 275773
rect 67465 275745 67499 275773
rect 67527 275745 67561 275773
rect 67589 275745 67623 275773
rect 67651 275745 67699 275773
rect 67389 266959 67699 275745
rect 67389 266931 67437 266959
rect 67465 266931 67499 266959
rect 67527 266931 67561 266959
rect 67589 266931 67623 266959
rect 67651 266931 67699 266959
rect 67389 266897 67699 266931
rect 67389 266869 67437 266897
rect 67465 266869 67499 266897
rect 67527 266869 67561 266897
rect 67589 266869 67623 266897
rect 67651 266869 67699 266897
rect 67389 266835 67699 266869
rect 67389 266807 67437 266835
rect 67465 266807 67499 266835
rect 67527 266807 67561 266835
rect 67589 266807 67623 266835
rect 67651 266807 67699 266835
rect 67389 266773 67699 266807
rect 67389 266745 67437 266773
rect 67465 266745 67499 266773
rect 67527 266745 67561 266773
rect 67589 266745 67623 266773
rect 67651 266745 67699 266773
rect 67389 257959 67699 266745
rect 67389 257931 67437 257959
rect 67465 257931 67499 257959
rect 67527 257931 67561 257959
rect 67589 257931 67623 257959
rect 67651 257931 67699 257959
rect 67389 257897 67699 257931
rect 67389 257869 67437 257897
rect 67465 257869 67499 257897
rect 67527 257869 67561 257897
rect 67589 257869 67623 257897
rect 67651 257869 67699 257897
rect 67389 257835 67699 257869
rect 67389 257807 67437 257835
rect 67465 257807 67499 257835
rect 67527 257807 67561 257835
rect 67589 257807 67623 257835
rect 67651 257807 67699 257835
rect 67389 257773 67699 257807
rect 67389 257745 67437 257773
rect 67465 257745 67499 257773
rect 67527 257745 67561 257773
rect 67589 257745 67623 257773
rect 67651 257745 67699 257773
rect 67389 254075 67699 257745
rect 74529 299190 74839 299718
rect 74529 299162 74577 299190
rect 74605 299162 74639 299190
rect 74667 299162 74701 299190
rect 74729 299162 74763 299190
rect 74791 299162 74839 299190
rect 74529 299128 74839 299162
rect 74529 299100 74577 299128
rect 74605 299100 74639 299128
rect 74667 299100 74701 299128
rect 74729 299100 74763 299128
rect 74791 299100 74839 299128
rect 74529 299066 74839 299100
rect 74529 299038 74577 299066
rect 74605 299038 74639 299066
rect 74667 299038 74701 299066
rect 74729 299038 74763 299066
rect 74791 299038 74839 299066
rect 74529 299004 74839 299038
rect 74529 298976 74577 299004
rect 74605 298976 74639 299004
rect 74667 298976 74701 299004
rect 74729 298976 74763 299004
rect 74791 298976 74839 299004
rect 74529 290959 74839 298976
rect 74529 290931 74577 290959
rect 74605 290931 74639 290959
rect 74667 290931 74701 290959
rect 74729 290931 74763 290959
rect 74791 290931 74839 290959
rect 74529 290897 74839 290931
rect 74529 290869 74577 290897
rect 74605 290869 74639 290897
rect 74667 290869 74701 290897
rect 74729 290869 74763 290897
rect 74791 290869 74839 290897
rect 74529 290835 74839 290869
rect 74529 290807 74577 290835
rect 74605 290807 74639 290835
rect 74667 290807 74701 290835
rect 74729 290807 74763 290835
rect 74791 290807 74839 290835
rect 74529 290773 74839 290807
rect 74529 290745 74577 290773
rect 74605 290745 74639 290773
rect 74667 290745 74701 290773
rect 74729 290745 74763 290773
rect 74791 290745 74839 290773
rect 74529 281959 74839 290745
rect 74529 281931 74577 281959
rect 74605 281931 74639 281959
rect 74667 281931 74701 281959
rect 74729 281931 74763 281959
rect 74791 281931 74839 281959
rect 74529 281897 74839 281931
rect 74529 281869 74577 281897
rect 74605 281869 74639 281897
rect 74667 281869 74701 281897
rect 74729 281869 74763 281897
rect 74791 281869 74839 281897
rect 74529 281835 74839 281869
rect 74529 281807 74577 281835
rect 74605 281807 74639 281835
rect 74667 281807 74701 281835
rect 74729 281807 74763 281835
rect 74791 281807 74839 281835
rect 74529 281773 74839 281807
rect 74529 281745 74577 281773
rect 74605 281745 74639 281773
rect 74667 281745 74701 281773
rect 74729 281745 74763 281773
rect 74791 281745 74839 281773
rect 74529 272959 74839 281745
rect 74529 272931 74577 272959
rect 74605 272931 74639 272959
rect 74667 272931 74701 272959
rect 74729 272931 74763 272959
rect 74791 272931 74839 272959
rect 74529 272897 74839 272931
rect 74529 272869 74577 272897
rect 74605 272869 74639 272897
rect 74667 272869 74701 272897
rect 74729 272869 74763 272897
rect 74791 272869 74839 272897
rect 74529 272835 74839 272869
rect 74529 272807 74577 272835
rect 74605 272807 74639 272835
rect 74667 272807 74701 272835
rect 74729 272807 74763 272835
rect 74791 272807 74839 272835
rect 74529 272773 74839 272807
rect 74529 272745 74577 272773
rect 74605 272745 74639 272773
rect 74667 272745 74701 272773
rect 74729 272745 74763 272773
rect 74791 272745 74839 272773
rect 74529 263959 74839 272745
rect 74529 263931 74577 263959
rect 74605 263931 74639 263959
rect 74667 263931 74701 263959
rect 74729 263931 74763 263959
rect 74791 263931 74839 263959
rect 74529 263897 74839 263931
rect 74529 263869 74577 263897
rect 74605 263869 74639 263897
rect 74667 263869 74701 263897
rect 74729 263869 74763 263897
rect 74791 263869 74839 263897
rect 74529 263835 74839 263869
rect 74529 263807 74577 263835
rect 74605 263807 74639 263835
rect 74667 263807 74701 263835
rect 74729 263807 74763 263835
rect 74791 263807 74839 263835
rect 74529 263773 74839 263807
rect 74529 263745 74577 263773
rect 74605 263745 74639 263773
rect 74667 263745 74701 263773
rect 74729 263745 74763 263773
rect 74791 263745 74839 263773
rect 74529 254959 74839 263745
rect 74529 254931 74577 254959
rect 74605 254931 74639 254959
rect 74667 254931 74701 254959
rect 74729 254931 74763 254959
rect 74791 254931 74839 254959
rect 74529 254897 74839 254931
rect 74529 254869 74577 254897
rect 74605 254869 74639 254897
rect 74667 254869 74701 254897
rect 74729 254869 74763 254897
rect 74791 254869 74839 254897
rect 74529 254835 74839 254869
rect 74529 254807 74577 254835
rect 74605 254807 74639 254835
rect 74667 254807 74701 254835
rect 74729 254807 74763 254835
rect 74791 254807 74839 254835
rect 74529 254773 74839 254807
rect 74529 254745 74577 254773
rect 74605 254745 74639 254773
rect 74667 254745 74701 254773
rect 74729 254745 74763 254773
rect 74791 254745 74839 254773
rect 74529 254075 74839 254745
rect 76389 299670 76699 299718
rect 76389 299642 76437 299670
rect 76465 299642 76499 299670
rect 76527 299642 76561 299670
rect 76589 299642 76623 299670
rect 76651 299642 76699 299670
rect 76389 299608 76699 299642
rect 76389 299580 76437 299608
rect 76465 299580 76499 299608
rect 76527 299580 76561 299608
rect 76589 299580 76623 299608
rect 76651 299580 76699 299608
rect 76389 299546 76699 299580
rect 76389 299518 76437 299546
rect 76465 299518 76499 299546
rect 76527 299518 76561 299546
rect 76589 299518 76623 299546
rect 76651 299518 76699 299546
rect 76389 299484 76699 299518
rect 76389 299456 76437 299484
rect 76465 299456 76499 299484
rect 76527 299456 76561 299484
rect 76589 299456 76623 299484
rect 76651 299456 76699 299484
rect 76389 293959 76699 299456
rect 76389 293931 76437 293959
rect 76465 293931 76499 293959
rect 76527 293931 76561 293959
rect 76589 293931 76623 293959
rect 76651 293931 76699 293959
rect 76389 293897 76699 293931
rect 76389 293869 76437 293897
rect 76465 293869 76499 293897
rect 76527 293869 76561 293897
rect 76589 293869 76623 293897
rect 76651 293869 76699 293897
rect 76389 293835 76699 293869
rect 76389 293807 76437 293835
rect 76465 293807 76499 293835
rect 76527 293807 76561 293835
rect 76589 293807 76623 293835
rect 76651 293807 76699 293835
rect 76389 293773 76699 293807
rect 76389 293745 76437 293773
rect 76465 293745 76499 293773
rect 76527 293745 76561 293773
rect 76589 293745 76623 293773
rect 76651 293745 76699 293773
rect 76389 284959 76699 293745
rect 76389 284931 76437 284959
rect 76465 284931 76499 284959
rect 76527 284931 76561 284959
rect 76589 284931 76623 284959
rect 76651 284931 76699 284959
rect 76389 284897 76699 284931
rect 76389 284869 76437 284897
rect 76465 284869 76499 284897
rect 76527 284869 76561 284897
rect 76589 284869 76623 284897
rect 76651 284869 76699 284897
rect 76389 284835 76699 284869
rect 76389 284807 76437 284835
rect 76465 284807 76499 284835
rect 76527 284807 76561 284835
rect 76589 284807 76623 284835
rect 76651 284807 76699 284835
rect 76389 284773 76699 284807
rect 76389 284745 76437 284773
rect 76465 284745 76499 284773
rect 76527 284745 76561 284773
rect 76589 284745 76623 284773
rect 76651 284745 76699 284773
rect 76389 275959 76699 284745
rect 76389 275931 76437 275959
rect 76465 275931 76499 275959
rect 76527 275931 76561 275959
rect 76589 275931 76623 275959
rect 76651 275931 76699 275959
rect 76389 275897 76699 275931
rect 76389 275869 76437 275897
rect 76465 275869 76499 275897
rect 76527 275869 76561 275897
rect 76589 275869 76623 275897
rect 76651 275869 76699 275897
rect 76389 275835 76699 275869
rect 76389 275807 76437 275835
rect 76465 275807 76499 275835
rect 76527 275807 76561 275835
rect 76589 275807 76623 275835
rect 76651 275807 76699 275835
rect 76389 275773 76699 275807
rect 76389 275745 76437 275773
rect 76465 275745 76499 275773
rect 76527 275745 76561 275773
rect 76589 275745 76623 275773
rect 76651 275745 76699 275773
rect 76389 266959 76699 275745
rect 76389 266931 76437 266959
rect 76465 266931 76499 266959
rect 76527 266931 76561 266959
rect 76589 266931 76623 266959
rect 76651 266931 76699 266959
rect 76389 266897 76699 266931
rect 76389 266869 76437 266897
rect 76465 266869 76499 266897
rect 76527 266869 76561 266897
rect 76589 266869 76623 266897
rect 76651 266869 76699 266897
rect 76389 266835 76699 266869
rect 76389 266807 76437 266835
rect 76465 266807 76499 266835
rect 76527 266807 76561 266835
rect 76589 266807 76623 266835
rect 76651 266807 76699 266835
rect 76389 266773 76699 266807
rect 76389 266745 76437 266773
rect 76465 266745 76499 266773
rect 76527 266745 76561 266773
rect 76589 266745 76623 266773
rect 76651 266745 76699 266773
rect 76389 257959 76699 266745
rect 76389 257931 76437 257959
rect 76465 257931 76499 257959
rect 76527 257931 76561 257959
rect 76589 257931 76623 257959
rect 76651 257931 76699 257959
rect 76389 257897 76699 257931
rect 76389 257869 76437 257897
rect 76465 257869 76499 257897
rect 76527 257869 76561 257897
rect 76589 257869 76623 257897
rect 76651 257869 76699 257897
rect 76389 257835 76699 257869
rect 76389 257807 76437 257835
rect 76465 257807 76499 257835
rect 76527 257807 76561 257835
rect 76589 257807 76623 257835
rect 76651 257807 76699 257835
rect 76389 257773 76699 257807
rect 76389 257745 76437 257773
rect 76465 257745 76499 257773
rect 76527 257745 76561 257773
rect 76589 257745 76623 257773
rect 76651 257745 76699 257773
rect 76389 254075 76699 257745
rect 83529 299190 83839 299718
rect 83529 299162 83577 299190
rect 83605 299162 83639 299190
rect 83667 299162 83701 299190
rect 83729 299162 83763 299190
rect 83791 299162 83839 299190
rect 83529 299128 83839 299162
rect 83529 299100 83577 299128
rect 83605 299100 83639 299128
rect 83667 299100 83701 299128
rect 83729 299100 83763 299128
rect 83791 299100 83839 299128
rect 83529 299066 83839 299100
rect 83529 299038 83577 299066
rect 83605 299038 83639 299066
rect 83667 299038 83701 299066
rect 83729 299038 83763 299066
rect 83791 299038 83839 299066
rect 83529 299004 83839 299038
rect 83529 298976 83577 299004
rect 83605 298976 83639 299004
rect 83667 298976 83701 299004
rect 83729 298976 83763 299004
rect 83791 298976 83839 299004
rect 83529 290959 83839 298976
rect 83529 290931 83577 290959
rect 83605 290931 83639 290959
rect 83667 290931 83701 290959
rect 83729 290931 83763 290959
rect 83791 290931 83839 290959
rect 83529 290897 83839 290931
rect 83529 290869 83577 290897
rect 83605 290869 83639 290897
rect 83667 290869 83701 290897
rect 83729 290869 83763 290897
rect 83791 290869 83839 290897
rect 83529 290835 83839 290869
rect 83529 290807 83577 290835
rect 83605 290807 83639 290835
rect 83667 290807 83701 290835
rect 83729 290807 83763 290835
rect 83791 290807 83839 290835
rect 83529 290773 83839 290807
rect 83529 290745 83577 290773
rect 83605 290745 83639 290773
rect 83667 290745 83701 290773
rect 83729 290745 83763 290773
rect 83791 290745 83839 290773
rect 83529 281959 83839 290745
rect 83529 281931 83577 281959
rect 83605 281931 83639 281959
rect 83667 281931 83701 281959
rect 83729 281931 83763 281959
rect 83791 281931 83839 281959
rect 83529 281897 83839 281931
rect 83529 281869 83577 281897
rect 83605 281869 83639 281897
rect 83667 281869 83701 281897
rect 83729 281869 83763 281897
rect 83791 281869 83839 281897
rect 83529 281835 83839 281869
rect 83529 281807 83577 281835
rect 83605 281807 83639 281835
rect 83667 281807 83701 281835
rect 83729 281807 83763 281835
rect 83791 281807 83839 281835
rect 83529 281773 83839 281807
rect 83529 281745 83577 281773
rect 83605 281745 83639 281773
rect 83667 281745 83701 281773
rect 83729 281745 83763 281773
rect 83791 281745 83839 281773
rect 83529 272959 83839 281745
rect 83529 272931 83577 272959
rect 83605 272931 83639 272959
rect 83667 272931 83701 272959
rect 83729 272931 83763 272959
rect 83791 272931 83839 272959
rect 83529 272897 83839 272931
rect 83529 272869 83577 272897
rect 83605 272869 83639 272897
rect 83667 272869 83701 272897
rect 83729 272869 83763 272897
rect 83791 272869 83839 272897
rect 83529 272835 83839 272869
rect 83529 272807 83577 272835
rect 83605 272807 83639 272835
rect 83667 272807 83701 272835
rect 83729 272807 83763 272835
rect 83791 272807 83839 272835
rect 83529 272773 83839 272807
rect 83529 272745 83577 272773
rect 83605 272745 83639 272773
rect 83667 272745 83701 272773
rect 83729 272745 83763 272773
rect 83791 272745 83839 272773
rect 83529 263959 83839 272745
rect 83529 263931 83577 263959
rect 83605 263931 83639 263959
rect 83667 263931 83701 263959
rect 83729 263931 83763 263959
rect 83791 263931 83839 263959
rect 83529 263897 83839 263931
rect 83529 263869 83577 263897
rect 83605 263869 83639 263897
rect 83667 263869 83701 263897
rect 83729 263869 83763 263897
rect 83791 263869 83839 263897
rect 83529 263835 83839 263869
rect 83529 263807 83577 263835
rect 83605 263807 83639 263835
rect 83667 263807 83701 263835
rect 83729 263807 83763 263835
rect 83791 263807 83839 263835
rect 83529 263773 83839 263807
rect 83529 263745 83577 263773
rect 83605 263745 83639 263773
rect 83667 263745 83701 263773
rect 83729 263745 83763 263773
rect 83791 263745 83839 263773
rect 83529 254959 83839 263745
rect 83529 254931 83577 254959
rect 83605 254931 83639 254959
rect 83667 254931 83701 254959
rect 83729 254931 83763 254959
rect 83791 254931 83839 254959
rect 83529 254897 83839 254931
rect 83529 254869 83577 254897
rect 83605 254869 83639 254897
rect 83667 254869 83701 254897
rect 83729 254869 83763 254897
rect 83791 254869 83839 254897
rect 83529 254835 83839 254869
rect 83529 254807 83577 254835
rect 83605 254807 83639 254835
rect 83667 254807 83701 254835
rect 83729 254807 83763 254835
rect 83791 254807 83839 254835
rect 83529 254773 83839 254807
rect 83529 254745 83577 254773
rect 83605 254745 83639 254773
rect 83667 254745 83701 254773
rect 83729 254745 83763 254773
rect 83791 254745 83839 254773
rect 83529 254075 83839 254745
rect 85389 299670 85699 299718
rect 85389 299642 85437 299670
rect 85465 299642 85499 299670
rect 85527 299642 85561 299670
rect 85589 299642 85623 299670
rect 85651 299642 85699 299670
rect 85389 299608 85699 299642
rect 85389 299580 85437 299608
rect 85465 299580 85499 299608
rect 85527 299580 85561 299608
rect 85589 299580 85623 299608
rect 85651 299580 85699 299608
rect 85389 299546 85699 299580
rect 85389 299518 85437 299546
rect 85465 299518 85499 299546
rect 85527 299518 85561 299546
rect 85589 299518 85623 299546
rect 85651 299518 85699 299546
rect 85389 299484 85699 299518
rect 85389 299456 85437 299484
rect 85465 299456 85499 299484
rect 85527 299456 85561 299484
rect 85589 299456 85623 299484
rect 85651 299456 85699 299484
rect 85389 293959 85699 299456
rect 85389 293931 85437 293959
rect 85465 293931 85499 293959
rect 85527 293931 85561 293959
rect 85589 293931 85623 293959
rect 85651 293931 85699 293959
rect 85389 293897 85699 293931
rect 85389 293869 85437 293897
rect 85465 293869 85499 293897
rect 85527 293869 85561 293897
rect 85589 293869 85623 293897
rect 85651 293869 85699 293897
rect 85389 293835 85699 293869
rect 85389 293807 85437 293835
rect 85465 293807 85499 293835
rect 85527 293807 85561 293835
rect 85589 293807 85623 293835
rect 85651 293807 85699 293835
rect 85389 293773 85699 293807
rect 85389 293745 85437 293773
rect 85465 293745 85499 293773
rect 85527 293745 85561 293773
rect 85589 293745 85623 293773
rect 85651 293745 85699 293773
rect 85389 284959 85699 293745
rect 85389 284931 85437 284959
rect 85465 284931 85499 284959
rect 85527 284931 85561 284959
rect 85589 284931 85623 284959
rect 85651 284931 85699 284959
rect 85389 284897 85699 284931
rect 85389 284869 85437 284897
rect 85465 284869 85499 284897
rect 85527 284869 85561 284897
rect 85589 284869 85623 284897
rect 85651 284869 85699 284897
rect 85389 284835 85699 284869
rect 85389 284807 85437 284835
rect 85465 284807 85499 284835
rect 85527 284807 85561 284835
rect 85589 284807 85623 284835
rect 85651 284807 85699 284835
rect 85389 284773 85699 284807
rect 85389 284745 85437 284773
rect 85465 284745 85499 284773
rect 85527 284745 85561 284773
rect 85589 284745 85623 284773
rect 85651 284745 85699 284773
rect 85389 275959 85699 284745
rect 85389 275931 85437 275959
rect 85465 275931 85499 275959
rect 85527 275931 85561 275959
rect 85589 275931 85623 275959
rect 85651 275931 85699 275959
rect 85389 275897 85699 275931
rect 85389 275869 85437 275897
rect 85465 275869 85499 275897
rect 85527 275869 85561 275897
rect 85589 275869 85623 275897
rect 85651 275869 85699 275897
rect 85389 275835 85699 275869
rect 85389 275807 85437 275835
rect 85465 275807 85499 275835
rect 85527 275807 85561 275835
rect 85589 275807 85623 275835
rect 85651 275807 85699 275835
rect 85389 275773 85699 275807
rect 85389 275745 85437 275773
rect 85465 275745 85499 275773
rect 85527 275745 85561 275773
rect 85589 275745 85623 275773
rect 85651 275745 85699 275773
rect 85389 266959 85699 275745
rect 85389 266931 85437 266959
rect 85465 266931 85499 266959
rect 85527 266931 85561 266959
rect 85589 266931 85623 266959
rect 85651 266931 85699 266959
rect 85389 266897 85699 266931
rect 85389 266869 85437 266897
rect 85465 266869 85499 266897
rect 85527 266869 85561 266897
rect 85589 266869 85623 266897
rect 85651 266869 85699 266897
rect 85389 266835 85699 266869
rect 85389 266807 85437 266835
rect 85465 266807 85499 266835
rect 85527 266807 85561 266835
rect 85589 266807 85623 266835
rect 85651 266807 85699 266835
rect 85389 266773 85699 266807
rect 85389 266745 85437 266773
rect 85465 266745 85499 266773
rect 85527 266745 85561 266773
rect 85589 266745 85623 266773
rect 85651 266745 85699 266773
rect 85389 257959 85699 266745
rect 85389 257931 85437 257959
rect 85465 257931 85499 257959
rect 85527 257931 85561 257959
rect 85589 257931 85623 257959
rect 85651 257931 85699 257959
rect 85389 257897 85699 257931
rect 85389 257869 85437 257897
rect 85465 257869 85499 257897
rect 85527 257869 85561 257897
rect 85589 257869 85623 257897
rect 85651 257869 85699 257897
rect 85389 257835 85699 257869
rect 85389 257807 85437 257835
rect 85465 257807 85499 257835
rect 85527 257807 85561 257835
rect 85589 257807 85623 257835
rect 85651 257807 85699 257835
rect 85389 257773 85699 257807
rect 85389 257745 85437 257773
rect 85465 257745 85499 257773
rect 85527 257745 85561 257773
rect 85589 257745 85623 257773
rect 85651 257745 85699 257773
rect 85389 254075 85699 257745
rect 92529 299190 92839 299718
rect 92529 299162 92577 299190
rect 92605 299162 92639 299190
rect 92667 299162 92701 299190
rect 92729 299162 92763 299190
rect 92791 299162 92839 299190
rect 92529 299128 92839 299162
rect 92529 299100 92577 299128
rect 92605 299100 92639 299128
rect 92667 299100 92701 299128
rect 92729 299100 92763 299128
rect 92791 299100 92839 299128
rect 92529 299066 92839 299100
rect 92529 299038 92577 299066
rect 92605 299038 92639 299066
rect 92667 299038 92701 299066
rect 92729 299038 92763 299066
rect 92791 299038 92839 299066
rect 92529 299004 92839 299038
rect 92529 298976 92577 299004
rect 92605 298976 92639 299004
rect 92667 298976 92701 299004
rect 92729 298976 92763 299004
rect 92791 298976 92839 299004
rect 92529 290959 92839 298976
rect 92529 290931 92577 290959
rect 92605 290931 92639 290959
rect 92667 290931 92701 290959
rect 92729 290931 92763 290959
rect 92791 290931 92839 290959
rect 92529 290897 92839 290931
rect 92529 290869 92577 290897
rect 92605 290869 92639 290897
rect 92667 290869 92701 290897
rect 92729 290869 92763 290897
rect 92791 290869 92839 290897
rect 92529 290835 92839 290869
rect 92529 290807 92577 290835
rect 92605 290807 92639 290835
rect 92667 290807 92701 290835
rect 92729 290807 92763 290835
rect 92791 290807 92839 290835
rect 92529 290773 92839 290807
rect 92529 290745 92577 290773
rect 92605 290745 92639 290773
rect 92667 290745 92701 290773
rect 92729 290745 92763 290773
rect 92791 290745 92839 290773
rect 92529 281959 92839 290745
rect 92529 281931 92577 281959
rect 92605 281931 92639 281959
rect 92667 281931 92701 281959
rect 92729 281931 92763 281959
rect 92791 281931 92839 281959
rect 92529 281897 92839 281931
rect 92529 281869 92577 281897
rect 92605 281869 92639 281897
rect 92667 281869 92701 281897
rect 92729 281869 92763 281897
rect 92791 281869 92839 281897
rect 92529 281835 92839 281869
rect 92529 281807 92577 281835
rect 92605 281807 92639 281835
rect 92667 281807 92701 281835
rect 92729 281807 92763 281835
rect 92791 281807 92839 281835
rect 92529 281773 92839 281807
rect 92529 281745 92577 281773
rect 92605 281745 92639 281773
rect 92667 281745 92701 281773
rect 92729 281745 92763 281773
rect 92791 281745 92839 281773
rect 92529 272959 92839 281745
rect 92529 272931 92577 272959
rect 92605 272931 92639 272959
rect 92667 272931 92701 272959
rect 92729 272931 92763 272959
rect 92791 272931 92839 272959
rect 92529 272897 92839 272931
rect 92529 272869 92577 272897
rect 92605 272869 92639 272897
rect 92667 272869 92701 272897
rect 92729 272869 92763 272897
rect 92791 272869 92839 272897
rect 92529 272835 92839 272869
rect 92529 272807 92577 272835
rect 92605 272807 92639 272835
rect 92667 272807 92701 272835
rect 92729 272807 92763 272835
rect 92791 272807 92839 272835
rect 92529 272773 92839 272807
rect 92529 272745 92577 272773
rect 92605 272745 92639 272773
rect 92667 272745 92701 272773
rect 92729 272745 92763 272773
rect 92791 272745 92839 272773
rect 92529 263959 92839 272745
rect 92529 263931 92577 263959
rect 92605 263931 92639 263959
rect 92667 263931 92701 263959
rect 92729 263931 92763 263959
rect 92791 263931 92839 263959
rect 92529 263897 92839 263931
rect 92529 263869 92577 263897
rect 92605 263869 92639 263897
rect 92667 263869 92701 263897
rect 92729 263869 92763 263897
rect 92791 263869 92839 263897
rect 92529 263835 92839 263869
rect 92529 263807 92577 263835
rect 92605 263807 92639 263835
rect 92667 263807 92701 263835
rect 92729 263807 92763 263835
rect 92791 263807 92839 263835
rect 92529 263773 92839 263807
rect 92529 263745 92577 263773
rect 92605 263745 92639 263773
rect 92667 263745 92701 263773
rect 92729 263745 92763 263773
rect 92791 263745 92839 263773
rect 92529 254959 92839 263745
rect 92529 254931 92577 254959
rect 92605 254931 92639 254959
rect 92667 254931 92701 254959
rect 92729 254931 92763 254959
rect 92791 254931 92839 254959
rect 92529 254897 92839 254931
rect 92529 254869 92577 254897
rect 92605 254869 92639 254897
rect 92667 254869 92701 254897
rect 92729 254869 92763 254897
rect 92791 254869 92839 254897
rect 92529 254835 92839 254869
rect 92529 254807 92577 254835
rect 92605 254807 92639 254835
rect 92667 254807 92701 254835
rect 92729 254807 92763 254835
rect 92791 254807 92839 254835
rect 92529 254773 92839 254807
rect 92529 254745 92577 254773
rect 92605 254745 92639 254773
rect 92667 254745 92701 254773
rect 92729 254745 92763 254773
rect 92791 254745 92839 254773
rect 92529 254075 92839 254745
rect 94389 299670 94699 299718
rect 94389 299642 94437 299670
rect 94465 299642 94499 299670
rect 94527 299642 94561 299670
rect 94589 299642 94623 299670
rect 94651 299642 94699 299670
rect 94389 299608 94699 299642
rect 94389 299580 94437 299608
rect 94465 299580 94499 299608
rect 94527 299580 94561 299608
rect 94589 299580 94623 299608
rect 94651 299580 94699 299608
rect 94389 299546 94699 299580
rect 94389 299518 94437 299546
rect 94465 299518 94499 299546
rect 94527 299518 94561 299546
rect 94589 299518 94623 299546
rect 94651 299518 94699 299546
rect 94389 299484 94699 299518
rect 94389 299456 94437 299484
rect 94465 299456 94499 299484
rect 94527 299456 94561 299484
rect 94589 299456 94623 299484
rect 94651 299456 94699 299484
rect 94389 293959 94699 299456
rect 94389 293931 94437 293959
rect 94465 293931 94499 293959
rect 94527 293931 94561 293959
rect 94589 293931 94623 293959
rect 94651 293931 94699 293959
rect 94389 293897 94699 293931
rect 94389 293869 94437 293897
rect 94465 293869 94499 293897
rect 94527 293869 94561 293897
rect 94589 293869 94623 293897
rect 94651 293869 94699 293897
rect 94389 293835 94699 293869
rect 94389 293807 94437 293835
rect 94465 293807 94499 293835
rect 94527 293807 94561 293835
rect 94589 293807 94623 293835
rect 94651 293807 94699 293835
rect 94389 293773 94699 293807
rect 94389 293745 94437 293773
rect 94465 293745 94499 293773
rect 94527 293745 94561 293773
rect 94589 293745 94623 293773
rect 94651 293745 94699 293773
rect 94389 284959 94699 293745
rect 94389 284931 94437 284959
rect 94465 284931 94499 284959
rect 94527 284931 94561 284959
rect 94589 284931 94623 284959
rect 94651 284931 94699 284959
rect 94389 284897 94699 284931
rect 94389 284869 94437 284897
rect 94465 284869 94499 284897
rect 94527 284869 94561 284897
rect 94589 284869 94623 284897
rect 94651 284869 94699 284897
rect 94389 284835 94699 284869
rect 94389 284807 94437 284835
rect 94465 284807 94499 284835
rect 94527 284807 94561 284835
rect 94589 284807 94623 284835
rect 94651 284807 94699 284835
rect 94389 284773 94699 284807
rect 94389 284745 94437 284773
rect 94465 284745 94499 284773
rect 94527 284745 94561 284773
rect 94589 284745 94623 284773
rect 94651 284745 94699 284773
rect 94389 275959 94699 284745
rect 94389 275931 94437 275959
rect 94465 275931 94499 275959
rect 94527 275931 94561 275959
rect 94589 275931 94623 275959
rect 94651 275931 94699 275959
rect 94389 275897 94699 275931
rect 94389 275869 94437 275897
rect 94465 275869 94499 275897
rect 94527 275869 94561 275897
rect 94589 275869 94623 275897
rect 94651 275869 94699 275897
rect 94389 275835 94699 275869
rect 94389 275807 94437 275835
rect 94465 275807 94499 275835
rect 94527 275807 94561 275835
rect 94589 275807 94623 275835
rect 94651 275807 94699 275835
rect 94389 275773 94699 275807
rect 94389 275745 94437 275773
rect 94465 275745 94499 275773
rect 94527 275745 94561 275773
rect 94589 275745 94623 275773
rect 94651 275745 94699 275773
rect 94389 266959 94699 275745
rect 94389 266931 94437 266959
rect 94465 266931 94499 266959
rect 94527 266931 94561 266959
rect 94589 266931 94623 266959
rect 94651 266931 94699 266959
rect 94389 266897 94699 266931
rect 94389 266869 94437 266897
rect 94465 266869 94499 266897
rect 94527 266869 94561 266897
rect 94589 266869 94623 266897
rect 94651 266869 94699 266897
rect 94389 266835 94699 266869
rect 94389 266807 94437 266835
rect 94465 266807 94499 266835
rect 94527 266807 94561 266835
rect 94589 266807 94623 266835
rect 94651 266807 94699 266835
rect 94389 266773 94699 266807
rect 94389 266745 94437 266773
rect 94465 266745 94499 266773
rect 94527 266745 94561 266773
rect 94589 266745 94623 266773
rect 94651 266745 94699 266773
rect 94389 257959 94699 266745
rect 94389 257931 94437 257959
rect 94465 257931 94499 257959
rect 94527 257931 94561 257959
rect 94589 257931 94623 257959
rect 94651 257931 94699 257959
rect 94389 257897 94699 257931
rect 94389 257869 94437 257897
rect 94465 257869 94499 257897
rect 94527 257869 94561 257897
rect 94589 257869 94623 257897
rect 94651 257869 94699 257897
rect 94389 257835 94699 257869
rect 94389 257807 94437 257835
rect 94465 257807 94499 257835
rect 94527 257807 94561 257835
rect 94589 257807 94623 257835
rect 94651 257807 94699 257835
rect 94389 257773 94699 257807
rect 94389 257745 94437 257773
rect 94465 257745 94499 257773
rect 94527 257745 94561 257773
rect 94589 257745 94623 257773
rect 94651 257745 94699 257773
rect 94389 254075 94699 257745
rect 101529 299190 101839 299718
rect 101529 299162 101577 299190
rect 101605 299162 101639 299190
rect 101667 299162 101701 299190
rect 101729 299162 101763 299190
rect 101791 299162 101839 299190
rect 101529 299128 101839 299162
rect 101529 299100 101577 299128
rect 101605 299100 101639 299128
rect 101667 299100 101701 299128
rect 101729 299100 101763 299128
rect 101791 299100 101839 299128
rect 101529 299066 101839 299100
rect 101529 299038 101577 299066
rect 101605 299038 101639 299066
rect 101667 299038 101701 299066
rect 101729 299038 101763 299066
rect 101791 299038 101839 299066
rect 101529 299004 101839 299038
rect 101529 298976 101577 299004
rect 101605 298976 101639 299004
rect 101667 298976 101701 299004
rect 101729 298976 101763 299004
rect 101791 298976 101839 299004
rect 101529 290959 101839 298976
rect 101529 290931 101577 290959
rect 101605 290931 101639 290959
rect 101667 290931 101701 290959
rect 101729 290931 101763 290959
rect 101791 290931 101839 290959
rect 101529 290897 101839 290931
rect 101529 290869 101577 290897
rect 101605 290869 101639 290897
rect 101667 290869 101701 290897
rect 101729 290869 101763 290897
rect 101791 290869 101839 290897
rect 101529 290835 101839 290869
rect 101529 290807 101577 290835
rect 101605 290807 101639 290835
rect 101667 290807 101701 290835
rect 101729 290807 101763 290835
rect 101791 290807 101839 290835
rect 101529 290773 101839 290807
rect 101529 290745 101577 290773
rect 101605 290745 101639 290773
rect 101667 290745 101701 290773
rect 101729 290745 101763 290773
rect 101791 290745 101839 290773
rect 101529 281959 101839 290745
rect 101529 281931 101577 281959
rect 101605 281931 101639 281959
rect 101667 281931 101701 281959
rect 101729 281931 101763 281959
rect 101791 281931 101839 281959
rect 101529 281897 101839 281931
rect 101529 281869 101577 281897
rect 101605 281869 101639 281897
rect 101667 281869 101701 281897
rect 101729 281869 101763 281897
rect 101791 281869 101839 281897
rect 101529 281835 101839 281869
rect 101529 281807 101577 281835
rect 101605 281807 101639 281835
rect 101667 281807 101701 281835
rect 101729 281807 101763 281835
rect 101791 281807 101839 281835
rect 101529 281773 101839 281807
rect 101529 281745 101577 281773
rect 101605 281745 101639 281773
rect 101667 281745 101701 281773
rect 101729 281745 101763 281773
rect 101791 281745 101839 281773
rect 101529 272959 101839 281745
rect 101529 272931 101577 272959
rect 101605 272931 101639 272959
rect 101667 272931 101701 272959
rect 101729 272931 101763 272959
rect 101791 272931 101839 272959
rect 101529 272897 101839 272931
rect 101529 272869 101577 272897
rect 101605 272869 101639 272897
rect 101667 272869 101701 272897
rect 101729 272869 101763 272897
rect 101791 272869 101839 272897
rect 101529 272835 101839 272869
rect 101529 272807 101577 272835
rect 101605 272807 101639 272835
rect 101667 272807 101701 272835
rect 101729 272807 101763 272835
rect 101791 272807 101839 272835
rect 101529 272773 101839 272807
rect 101529 272745 101577 272773
rect 101605 272745 101639 272773
rect 101667 272745 101701 272773
rect 101729 272745 101763 272773
rect 101791 272745 101839 272773
rect 101529 263959 101839 272745
rect 101529 263931 101577 263959
rect 101605 263931 101639 263959
rect 101667 263931 101701 263959
rect 101729 263931 101763 263959
rect 101791 263931 101839 263959
rect 101529 263897 101839 263931
rect 101529 263869 101577 263897
rect 101605 263869 101639 263897
rect 101667 263869 101701 263897
rect 101729 263869 101763 263897
rect 101791 263869 101839 263897
rect 101529 263835 101839 263869
rect 101529 263807 101577 263835
rect 101605 263807 101639 263835
rect 101667 263807 101701 263835
rect 101729 263807 101763 263835
rect 101791 263807 101839 263835
rect 101529 263773 101839 263807
rect 101529 263745 101577 263773
rect 101605 263745 101639 263773
rect 101667 263745 101701 263773
rect 101729 263745 101763 263773
rect 101791 263745 101839 263773
rect 101529 254959 101839 263745
rect 101529 254931 101577 254959
rect 101605 254931 101639 254959
rect 101667 254931 101701 254959
rect 101729 254931 101763 254959
rect 101791 254931 101839 254959
rect 101529 254897 101839 254931
rect 101529 254869 101577 254897
rect 101605 254869 101639 254897
rect 101667 254869 101701 254897
rect 101729 254869 101763 254897
rect 101791 254869 101839 254897
rect 101529 254835 101839 254869
rect 101529 254807 101577 254835
rect 101605 254807 101639 254835
rect 101667 254807 101701 254835
rect 101729 254807 101763 254835
rect 101791 254807 101839 254835
rect 101529 254773 101839 254807
rect 101529 254745 101577 254773
rect 101605 254745 101639 254773
rect 101667 254745 101701 254773
rect 101729 254745 101763 254773
rect 101791 254745 101839 254773
rect 101529 254394 101839 254745
rect 103389 299670 103699 299718
rect 103389 299642 103437 299670
rect 103465 299642 103499 299670
rect 103527 299642 103561 299670
rect 103589 299642 103623 299670
rect 103651 299642 103699 299670
rect 103389 299608 103699 299642
rect 103389 299580 103437 299608
rect 103465 299580 103499 299608
rect 103527 299580 103561 299608
rect 103589 299580 103623 299608
rect 103651 299580 103699 299608
rect 103389 299546 103699 299580
rect 103389 299518 103437 299546
rect 103465 299518 103499 299546
rect 103527 299518 103561 299546
rect 103589 299518 103623 299546
rect 103651 299518 103699 299546
rect 103389 299484 103699 299518
rect 103389 299456 103437 299484
rect 103465 299456 103499 299484
rect 103527 299456 103561 299484
rect 103589 299456 103623 299484
rect 103651 299456 103699 299484
rect 103389 293959 103699 299456
rect 103389 293931 103437 293959
rect 103465 293931 103499 293959
rect 103527 293931 103561 293959
rect 103589 293931 103623 293959
rect 103651 293931 103699 293959
rect 103389 293897 103699 293931
rect 103389 293869 103437 293897
rect 103465 293869 103499 293897
rect 103527 293869 103561 293897
rect 103589 293869 103623 293897
rect 103651 293869 103699 293897
rect 103389 293835 103699 293869
rect 103389 293807 103437 293835
rect 103465 293807 103499 293835
rect 103527 293807 103561 293835
rect 103589 293807 103623 293835
rect 103651 293807 103699 293835
rect 103389 293773 103699 293807
rect 103389 293745 103437 293773
rect 103465 293745 103499 293773
rect 103527 293745 103561 293773
rect 103589 293745 103623 293773
rect 103651 293745 103699 293773
rect 103389 284959 103699 293745
rect 103389 284931 103437 284959
rect 103465 284931 103499 284959
rect 103527 284931 103561 284959
rect 103589 284931 103623 284959
rect 103651 284931 103699 284959
rect 103389 284897 103699 284931
rect 103389 284869 103437 284897
rect 103465 284869 103499 284897
rect 103527 284869 103561 284897
rect 103589 284869 103623 284897
rect 103651 284869 103699 284897
rect 103389 284835 103699 284869
rect 103389 284807 103437 284835
rect 103465 284807 103499 284835
rect 103527 284807 103561 284835
rect 103589 284807 103623 284835
rect 103651 284807 103699 284835
rect 103389 284773 103699 284807
rect 103389 284745 103437 284773
rect 103465 284745 103499 284773
rect 103527 284745 103561 284773
rect 103589 284745 103623 284773
rect 103651 284745 103699 284773
rect 103389 275959 103699 284745
rect 103389 275931 103437 275959
rect 103465 275931 103499 275959
rect 103527 275931 103561 275959
rect 103589 275931 103623 275959
rect 103651 275931 103699 275959
rect 103389 275897 103699 275931
rect 103389 275869 103437 275897
rect 103465 275869 103499 275897
rect 103527 275869 103561 275897
rect 103589 275869 103623 275897
rect 103651 275869 103699 275897
rect 103389 275835 103699 275869
rect 103389 275807 103437 275835
rect 103465 275807 103499 275835
rect 103527 275807 103561 275835
rect 103589 275807 103623 275835
rect 103651 275807 103699 275835
rect 103389 275773 103699 275807
rect 103389 275745 103437 275773
rect 103465 275745 103499 275773
rect 103527 275745 103561 275773
rect 103589 275745 103623 275773
rect 103651 275745 103699 275773
rect 103389 266959 103699 275745
rect 103389 266931 103437 266959
rect 103465 266931 103499 266959
rect 103527 266931 103561 266959
rect 103589 266931 103623 266959
rect 103651 266931 103699 266959
rect 103389 266897 103699 266931
rect 103389 266869 103437 266897
rect 103465 266869 103499 266897
rect 103527 266869 103561 266897
rect 103589 266869 103623 266897
rect 103651 266869 103699 266897
rect 103389 266835 103699 266869
rect 103389 266807 103437 266835
rect 103465 266807 103499 266835
rect 103527 266807 103561 266835
rect 103589 266807 103623 266835
rect 103651 266807 103699 266835
rect 103389 266773 103699 266807
rect 103389 266745 103437 266773
rect 103465 266745 103499 266773
rect 103527 266745 103561 266773
rect 103589 266745 103623 266773
rect 103651 266745 103699 266773
rect 103389 257959 103699 266745
rect 103389 257931 103437 257959
rect 103465 257931 103499 257959
rect 103527 257931 103561 257959
rect 103589 257931 103623 257959
rect 103651 257931 103699 257959
rect 103389 257897 103699 257931
rect 103389 257869 103437 257897
rect 103465 257869 103499 257897
rect 103527 257869 103561 257897
rect 103589 257869 103623 257897
rect 103651 257869 103699 257897
rect 103389 257835 103699 257869
rect 103389 257807 103437 257835
rect 103465 257807 103499 257835
rect 103527 257807 103561 257835
rect 103589 257807 103623 257835
rect 103651 257807 103699 257835
rect 103389 257773 103699 257807
rect 103389 257745 103437 257773
rect 103465 257745 103499 257773
rect 103527 257745 103561 257773
rect 103589 257745 103623 257773
rect 103651 257745 103699 257773
rect 103389 254075 103699 257745
rect 110529 299190 110839 299718
rect 110529 299162 110577 299190
rect 110605 299162 110639 299190
rect 110667 299162 110701 299190
rect 110729 299162 110763 299190
rect 110791 299162 110839 299190
rect 110529 299128 110839 299162
rect 110529 299100 110577 299128
rect 110605 299100 110639 299128
rect 110667 299100 110701 299128
rect 110729 299100 110763 299128
rect 110791 299100 110839 299128
rect 110529 299066 110839 299100
rect 110529 299038 110577 299066
rect 110605 299038 110639 299066
rect 110667 299038 110701 299066
rect 110729 299038 110763 299066
rect 110791 299038 110839 299066
rect 110529 299004 110839 299038
rect 110529 298976 110577 299004
rect 110605 298976 110639 299004
rect 110667 298976 110701 299004
rect 110729 298976 110763 299004
rect 110791 298976 110839 299004
rect 110529 290959 110839 298976
rect 110529 290931 110577 290959
rect 110605 290931 110639 290959
rect 110667 290931 110701 290959
rect 110729 290931 110763 290959
rect 110791 290931 110839 290959
rect 110529 290897 110839 290931
rect 110529 290869 110577 290897
rect 110605 290869 110639 290897
rect 110667 290869 110701 290897
rect 110729 290869 110763 290897
rect 110791 290869 110839 290897
rect 110529 290835 110839 290869
rect 110529 290807 110577 290835
rect 110605 290807 110639 290835
rect 110667 290807 110701 290835
rect 110729 290807 110763 290835
rect 110791 290807 110839 290835
rect 110529 290773 110839 290807
rect 110529 290745 110577 290773
rect 110605 290745 110639 290773
rect 110667 290745 110701 290773
rect 110729 290745 110763 290773
rect 110791 290745 110839 290773
rect 110529 281959 110839 290745
rect 110529 281931 110577 281959
rect 110605 281931 110639 281959
rect 110667 281931 110701 281959
rect 110729 281931 110763 281959
rect 110791 281931 110839 281959
rect 110529 281897 110839 281931
rect 110529 281869 110577 281897
rect 110605 281869 110639 281897
rect 110667 281869 110701 281897
rect 110729 281869 110763 281897
rect 110791 281869 110839 281897
rect 110529 281835 110839 281869
rect 110529 281807 110577 281835
rect 110605 281807 110639 281835
rect 110667 281807 110701 281835
rect 110729 281807 110763 281835
rect 110791 281807 110839 281835
rect 110529 281773 110839 281807
rect 110529 281745 110577 281773
rect 110605 281745 110639 281773
rect 110667 281745 110701 281773
rect 110729 281745 110763 281773
rect 110791 281745 110839 281773
rect 110529 272959 110839 281745
rect 110529 272931 110577 272959
rect 110605 272931 110639 272959
rect 110667 272931 110701 272959
rect 110729 272931 110763 272959
rect 110791 272931 110839 272959
rect 110529 272897 110839 272931
rect 110529 272869 110577 272897
rect 110605 272869 110639 272897
rect 110667 272869 110701 272897
rect 110729 272869 110763 272897
rect 110791 272869 110839 272897
rect 110529 272835 110839 272869
rect 110529 272807 110577 272835
rect 110605 272807 110639 272835
rect 110667 272807 110701 272835
rect 110729 272807 110763 272835
rect 110791 272807 110839 272835
rect 110529 272773 110839 272807
rect 110529 272745 110577 272773
rect 110605 272745 110639 272773
rect 110667 272745 110701 272773
rect 110729 272745 110763 272773
rect 110791 272745 110839 272773
rect 110529 263959 110839 272745
rect 110529 263931 110577 263959
rect 110605 263931 110639 263959
rect 110667 263931 110701 263959
rect 110729 263931 110763 263959
rect 110791 263931 110839 263959
rect 110529 263897 110839 263931
rect 110529 263869 110577 263897
rect 110605 263869 110639 263897
rect 110667 263869 110701 263897
rect 110729 263869 110763 263897
rect 110791 263869 110839 263897
rect 110529 263835 110839 263869
rect 110529 263807 110577 263835
rect 110605 263807 110639 263835
rect 110667 263807 110701 263835
rect 110729 263807 110763 263835
rect 110791 263807 110839 263835
rect 110529 263773 110839 263807
rect 110529 263745 110577 263773
rect 110605 263745 110639 263773
rect 110667 263745 110701 263773
rect 110729 263745 110763 263773
rect 110791 263745 110839 263773
rect 110529 254959 110839 263745
rect 110529 254931 110577 254959
rect 110605 254931 110639 254959
rect 110667 254931 110701 254959
rect 110729 254931 110763 254959
rect 110791 254931 110839 254959
rect 110529 254897 110839 254931
rect 110529 254869 110577 254897
rect 110605 254869 110639 254897
rect 110667 254869 110701 254897
rect 110729 254869 110763 254897
rect 110791 254869 110839 254897
rect 110529 254835 110839 254869
rect 110529 254807 110577 254835
rect 110605 254807 110639 254835
rect 110667 254807 110701 254835
rect 110729 254807 110763 254835
rect 110791 254807 110839 254835
rect 110529 254773 110839 254807
rect 110529 254745 110577 254773
rect 110605 254745 110639 254773
rect 110667 254745 110701 254773
rect 110729 254745 110763 254773
rect 110791 254745 110839 254773
rect 110529 254075 110839 254745
rect 112389 299670 112699 299718
rect 112389 299642 112437 299670
rect 112465 299642 112499 299670
rect 112527 299642 112561 299670
rect 112589 299642 112623 299670
rect 112651 299642 112699 299670
rect 112389 299608 112699 299642
rect 112389 299580 112437 299608
rect 112465 299580 112499 299608
rect 112527 299580 112561 299608
rect 112589 299580 112623 299608
rect 112651 299580 112699 299608
rect 112389 299546 112699 299580
rect 112389 299518 112437 299546
rect 112465 299518 112499 299546
rect 112527 299518 112561 299546
rect 112589 299518 112623 299546
rect 112651 299518 112699 299546
rect 112389 299484 112699 299518
rect 112389 299456 112437 299484
rect 112465 299456 112499 299484
rect 112527 299456 112561 299484
rect 112589 299456 112623 299484
rect 112651 299456 112699 299484
rect 112389 293959 112699 299456
rect 112389 293931 112437 293959
rect 112465 293931 112499 293959
rect 112527 293931 112561 293959
rect 112589 293931 112623 293959
rect 112651 293931 112699 293959
rect 112389 293897 112699 293931
rect 112389 293869 112437 293897
rect 112465 293869 112499 293897
rect 112527 293869 112561 293897
rect 112589 293869 112623 293897
rect 112651 293869 112699 293897
rect 112389 293835 112699 293869
rect 112389 293807 112437 293835
rect 112465 293807 112499 293835
rect 112527 293807 112561 293835
rect 112589 293807 112623 293835
rect 112651 293807 112699 293835
rect 112389 293773 112699 293807
rect 112389 293745 112437 293773
rect 112465 293745 112499 293773
rect 112527 293745 112561 293773
rect 112589 293745 112623 293773
rect 112651 293745 112699 293773
rect 112389 284959 112699 293745
rect 112389 284931 112437 284959
rect 112465 284931 112499 284959
rect 112527 284931 112561 284959
rect 112589 284931 112623 284959
rect 112651 284931 112699 284959
rect 112389 284897 112699 284931
rect 112389 284869 112437 284897
rect 112465 284869 112499 284897
rect 112527 284869 112561 284897
rect 112589 284869 112623 284897
rect 112651 284869 112699 284897
rect 112389 284835 112699 284869
rect 112389 284807 112437 284835
rect 112465 284807 112499 284835
rect 112527 284807 112561 284835
rect 112589 284807 112623 284835
rect 112651 284807 112699 284835
rect 112389 284773 112699 284807
rect 112389 284745 112437 284773
rect 112465 284745 112499 284773
rect 112527 284745 112561 284773
rect 112589 284745 112623 284773
rect 112651 284745 112699 284773
rect 112389 275959 112699 284745
rect 112389 275931 112437 275959
rect 112465 275931 112499 275959
rect 112527 275931 112561 275959
rect 112589 275931 112623 275959
rect 112651 275931 112699 275959
rect 112389 275897 112699 275931
rect 112389 275869 112437 275897
rect 112465 275869 112499 275897
rect 112527 275869 112561 275897
rect 112589 275869 112623 275897
rect 112651 275869 112699 275897
rect 112389 275835 112699 275869
rect 112389 275807 112437 275835
rect 112465 275807 112499 275835
rect 112527 275807 112561 275835
rect 112589 275807 112623 275835
rect 112651 275807 112699 275835
rect 112389 275773 112699 275807
rect 112389 275745 112437 275773
rect 112465 275745 112499 275773
rect 112527 275745 112561 275773
rect 112589 275745 112623 275773
rect 112651 275745 112699 275773
rect 112389 266959 112699 275745
rect 112389 266931 112437 266959
rect 112465 266931 112499 266959
rect 112527 266931 112561 266959
rect 112589 266931 112623 266959
rect 112651 266931 112699 266959
rect 112389 266897 112699 266931
rect 112389 266869 112437 266897
rect 112465 266869 112499 266897
rect 112527 266869 112561 266897
rect 112589 266869 112623 266897
rect 112651 266869 112699 266897
rect 112389 266835 112699 266869
rect 112389 266807 112437 266835
rect 112465 266807 112499 266835
rect 112527 266807 112561 266835
rect 112589 266807 112623 266835
rect 112651 266807 112699 266835
rect 112389 266773 112699 266807
rect 112389 266745 112437 266773
rect 112465 266745 112499 266773
rect 112527 266745 112561 266773
rect 112589 266745 112623 266773
rect 112651 266745 112699 266773
rect 112389 257959 112699 266745
rect 112389 257931 112437 257959
rect 112465 257931 112499 257959
rect 112527 257931 112561 257959
rect 112589 257931 112623 257959
rect 112651 257931 112699 257959
rect 112389 257897 112699 257931
rect 112389 257869 112437 257897
rect 112465 257869 112499 257897
rect 112527 257869 112561 257897
rect 112589 257869 112623 257897
rect 112651 257869 112699 257897
rect 112389 257835 112699 257869
rect 112389 257807 112437 257835
rect 112465 257807 112499 257835
rect 112527 257807 112561 257835
rect 112589 257807 112623 257835
rect 112651 257807 112699 257835
rect 112389 257773 112699 257807
rect 112389 257745 112437 257773
rect 112465 257745 112499 257773
rect 112527 257745 112561 257773
rect 112589 257745 112623 257773
rect 112651 257745 112699 257773
rect 112389 254075 112699 257745
rect 119529 299190 119839 299718
rect 119529 299162 119577 299190
rect 119605 299162 119639 299190
rect 119667 299162 119701 299190
rect 119729 299162 119763 299190
rect 119791 299162 119839 299190
rect 119529 299128 119839 299162
rect 119529 299100 119577 299128
rect 119605 299100 119639 299128
rect 119667 299100 119701 299128
rect 119729 299100 119763 299128
rect 119791 299100 119839 299128
rect 119529 299066 119839 299100
rect 119529 299038 119577 299066
rect 119605 299038 119639 299066
rect 119667 299038 119701 299066
rect 119729 299038 119763 299066
rect 119791 299038 119839 299066
rect 119529 299004 119839 299038
rect 119529 298976 119577 299004
rect 119605 298976 119639 299004
rect 119667 298976 119701 299004
rect 119729 298976 119763 299004
rect 119791 298976 119839 299004
rect 119529 290959 119839 298976
rect 119529 290931 119577 290959
rect 119605 290931 119639 290959
rect 119667 290931 119701 290959
rect 119729 290931 119763 290959
rect 119791 290931 119839 290959
rect 119529 290897 119839 290931
rect 119529 290869 119577 290897
rect 119605 290869 119639 290897
rect 119667 290869 119701 290897
rect 119729 290869 119763 290897
rect 119791 290869 119839 290897
rect 119529 290835 119839 290869
rect 119529 290807 119577 290835
rect 119605 290807 119639 290835
rect 119667 290807 119701 290835
rect 119729 290807 119763 290835
rect 119791 290807 119839 290835
rect 119529 290773 119839 290807
rect 119529 290745 119577 290773
rect 119605 290745 119639 290773
rect 119667 290745 119701 290773
rect 119729 290745 119763 290773
rect 119791 290745 119839 290773
rect 119529 281959 119839 290745
rect 119529 281931 119577 281959
rect 119605 281931 119639 281959
rect 119667 281931 119701 281959
rect 119729 281931 119763 281959
rect 119791 281931 119839 281959
rect 119529 281897 119839 281931
rect 119529 281869 119577 281897
rect 119605 281869 119639 281897
rect 119667 281869 119701 281897
rect 119729 281869 119763 281897
rect 119791 281869 119839 281897
rect 119529 281835 119839 281869
rect 119529 281807 119577 281835
rect 119605 281807 119639 281835
rect 119667 281807 119701 281835
rect 119729 281807 119763 281835
rect 119791 281807 119839 281835
rect 119529 281773 119839 281807
rect 119529 281745 119577 281773
rect 119605 281745 119639 281773
rect 119667 281745 119701 281773
rect 119729 281745 119763 281773
rect 119791 281745 119839 281773
rect 119529 272959 119839 281745
rect 119529 272931 119577 272959
rect 119605 272931 119639 272959
rect 119667 272931 119701 272959
rect 119729 272931 119763 272959
rect 119791 272931 119839 272959
rect 119529 272897 119839 272931
rect 119529 272869 119577 272897
rect 119605 272869 119639 272897
rect 119667 272869 119701 272897
rect 119729 272869 119763 272897
rect 119791 272869 119839 272897
rect 119529 272835 119839 272869
rect 119529 272807 119577 272835
rect 119605 272807 119639 272835
rect 119667 272807 119701 272835
rect 119729 272807 119763 272835
rect 119791 272807 119839 272835
rect 119529 272773 119839 272807
rect 119529 272745 119577 272773
rect 119605 272745 119639 272773
rect 119667 272745 119701 272773
rect 119729 272745 119763 272773
rect 119791 272745 119839 272773
rect 119529 263959 119839 272745
rect 119529 263931 119577 263959
rect 119605 263931 119639 263959
rect 119667 263931 119701 263959
rect 119729 263931 119763 263959
rect 119791 263931 119839 263959
rect 119529 263897 119839 263931
rect 119529 263869 119577 263897
rect 119605 263869 119639 263897
rect 119667 263869 119701 263897
rect 119729 263869 119763 263897
rect 119791 263869 119839 263897
rect 119529 263835 119839 263869
rect 119529 263807 119577 263835
rect 119605 263807 119639 263835
rect 119667 263807 119701 263835
rect 119729 263807 119763 263835
rect 119791 263807 119839 263835
rect 119529 263773 119839 263807
rect 119529 263745 119577 263773
rect 119605 263745 119639 263773
rect 119667 263745 119701 263773
rect 119729 263745 119763 263773
rect 119791 263745 119839 263773
rect 119529 254959 119839 263745
rect 119529 254931 119577 254959
rect 119605 254931 119639 254959
rect 119667 254931 119701 254959
rect 119729 254931 119763 254959
rect 119791 254931 119839 254959
rect 119529 254897 119839 254931
rect 119529 254869 119577 254897
rect 119605 254869 119639 254897
rect 119667 254869 119701 254897
rect 119729 254869 119763 254897
rect 119791 254869 119839 254897
rect 119529 254835 119839 254869
rect 119529 254807 119577 254835
rect 119605 254807 119639 254835
rect 119667 254807 119701 254835
rect 119729 254807 119763 254835
rect 119791 254807 119839 254835
rect 119529 254773 119839 254807
rect 119529 254745 119577 254773
rect 119605 254745 119639 254773
rect 119667 254745 119701 254773
rect 119729 254745 119763 254773
rect 119791 254745 119839 254773
rect 119529 254075 119839 254745
rect 121389 299670 121699 299718
rect 121389 299642 121437 299670
rect 121465 299642 121499 299670
rect 121527 299642 121561 299670
rect 121589 299642 121623 299670
rect 121651 299642 121699 299670
rect 121389 299608 121699 299642
rect 121389 299580 121437 299608
rect 121465 299580 121499 299608
rect 121527 299580 121561 299608
rect 121589 299580 121623 299608
rect 121651 299580 121699 299608
rect 121389 299546 121699 299580
rect 121389 299518 121437 299546
rect 121465 299518 121499 299546
rect 121527 299518 121561 299546
rect 121589 299518 121623 299546
rect 121651 299518 121699 299546
rect 121389 299484 121699 299518
rect 121389 299456 121437 299484
rect 121465 299456 121499 299484
rect 121527 299456 121561 299484
rect 121589 299456 121623 299484
rect 121651 299456 121699 299484
rect 121389 293959 121699 299456
rect 121389 293931 121437 293959
rect 121465 293931 121499 293959
rect 121527 293931 121561 293959
rect 121589 293931 121623 293959
rect 121651 293931 121699 293959
rect 121389 293897 121699 293931
rect 121389 293869 121437 293897
rect 121465 293869 121499 293897
rect 121527 293869 121561 293897
rect 121589 293869 121623 293897
rect 121651 293869 121699 293897
rect 121389 293835 121699 293869
rect 121389 293807 121437 293835
rect 121465 293807 121499 293835
rect 121527 293807 121561 293835
rect 121589 293807 121623 293835
rect 121651 293807 121699 293835
rect 121389 293773 121699 293807
rect 121389 293745 121437 293773
rect 121465 293745 121499 293773
rect 121527 293745 121561 293773
rect 121589 293745 121623 293773
rect 121651 293745 121699 293773
rect 121389 284959 121699 293745
rect 121389 284931 121437 284959
rect 121465 284931 121499 284959
rect 121527 284931 121561 284959
rect 121589 284931 121623 284959
rect 121651 284931 121699 284959
rect 121389 284897 121699 284931
rect 121389 284869 121437 284897
rect 121465 284869 121499 284897
rect 121527 284869 121561 284897
rect 121589 284869 121623 284897
rect 121651 284869 121699 284897
rect 121389 284835 121699 284869
rect 121389 284807 121437 284835
rect 121465 284807 121499 284835
rect 121527 284807 121561 284835
rect 121589 284807 121623 284835
rect 121651 284807 121699 284835
rect 121389 284773 121699 284807
rect 121389 284745 121437 284773
rect 121465 284745 121499 284773
rect 121527 284745 121561 284773
rect 121589 284745 121623 284773
rect 121651 284745 121699 284773
rect 121389 275959 121699 284745
rect 121389 275931 121437 275959
rect 121465 275931 121499 275959
rect 121527 275931 121561 275959
rect 121589 275931 121623 275959
rect 121651 275931 121699 275959
rect 121389 275897 121699 275931
rect 121389 275869 121437 275897
rect 121465 275869 121499 275897
rect 121527 275869 121561 275897
rect 121589 275869 121623 275897
rect 121651 275869 121699 275897
rect 121389 275835 121699 275869
rect 121389 275807 121437 275835
rect 121465 275807 121499 275835
rect 121527 275807 121561 275835
rect 121589 275807 121623 275835
rect 121651 275807 121699 275835
rect 121389 275773 121699 275807
rect 121389 275745 121437 275773
rect 121465 275745 121499 275773
rect 121527 275745 121561 275773
rect 121589 275745 121623 275773
rect 121651 275745 121699 275773
rect 121389 266959 121699 275745
rect 121389 266931 121437 266959
rect 121465 266931 121499 266959
rect 121527 266931 121561 266959
rect 121589 266931 121623 266959
rect 121651 266931 121699 266959
rect 121389 266897 121699 266931
rect 121389 266869 121437 266897
rect 121465 266869 121499 266897
rect 121527 266869 121561 266897
rect 121589 266869 121623 266897
rect 121651 266869 121699 266897
rect 121389 266835 121699 266869
rect 121389 266807 121437 266835
rect 121465 266807 121499 266835
rect 121527 266807 121561 266835
rect 121589 266807 121623 266835
rect 121651 266807 121699 266835
rect 121389 266773 121699 266807
rect 121389 266745 121437 266773
rect 121465 266745 121499 266773
rect 121527 266745 121561 266773
rect 121589 266745 121623 266773
rect 121651 266745 121699 266773
rect 121389 257959 121699 266745
rect 121389 257931 121437 257959
rect 121465 257931 121499 257959
rect 121527 257931 121561 257959
rect 121589 257931 121623 257959
rect 121651 257931 121699 257959
rect 121389 257897 121699 257931
rect 121389 257869 121437 257897
rect 121465 257869 121499 257897
rect 121527 257869 121561 257897
rect 121589 257869 121623 257897
rect 121651 257869 121699 257897
rect 121389 257835 121699 257869
rect 121389 257807 121437 257835
rect 121465 257807 121499 257835
rect 121527 257807 121561 257835
rect 121589 257807 121623 257835
rect 121651 257807 121699 257835
rect 121389 257773 121699 257807
rect 121389 257745 121437 257773
rect 121465 257745 121499 257773
rect 121527 257745 121561 257773
rect 121589 257745 121623 257773
rect 121651 257745 121699 257773
rect 121389 254075 121699 257745
rect 128529 299190 128839 299718
rect 128529 299162 128577 299190
rect 128605 299162 128639 299190
rect 128667 299162 128701 299190
rect 128729 299162 128763 299190
rect 128791 299162 128839 299190
rect 128529 299128 128839 299162
rect 128529 299100 128577 299128
rect 128605 299100 128639 299128
rect 128667 299100 128701 299128
rect 128729 299100 128763 299128
rect 128791 299100 128839 299128
rect 128529 299066 128839 299100
rect 128529 299038 128577 299066
rect 128605 299038 128639 299066
rect 128667 299038 128701 299066
rect 128729 299038 128763 299066
rect 128791 299038 128839 299066
rect 128529 299004 128839 299038
rect 128529 298976 128577 299004
rect 128605 298976 128639 299004
rect 128667 298976 128701 299004
rect 128729 298976 128763 299004
rect 128791 298976 128839 299004
rect 128529 290959 128839 298976
rect 128529 290931 128577 290959
rect 128605 290931 128639 290959
rect 128667 290931 128701 290959
rect 128729 290931 128763 290959
rect 128791 290931 128839 290959
rect 128529 290897 128839 290931
rect 128529 290869 128577 290897
rect 128605 290869 128639 290897
rect 128667 290869 128701 290897
rect 128729 290869 128763 290897
rect 128791 290869 128839 290897
rect 128529 290835 128839 290869
rect 128529 290807 128577 290835
rect 128605 290807 128639 290835
rect 128667 290807 128701 290835
rect 128729 290807 128763 290835
rect 128791 290807 128839 290835
rect 128529 290773 128839 290807
rect 128529 290745 128577 290773
rect 128605 290745 128639 290773
rect 128667 290745 128701 290773
rect 128729 290745 128763 290773
rect 128791 290745 128839 290773
rect 128529 281959 128839 290745
rect 128529 281931 128577 281959
rect 128605 281931 128639 281959
rect 128667 281931 128701 281959
rect 128729 281931 128763 281959
rect 128791 281931 128839 281959
rect 128529 281897 128839 281931
rect 128529 281869 128577 281897
rect 128605 281869 128639 281897
rect 128667 281869 128701 281897
rect 128729 281869 128763 281897
rect 128791 281869 128839 281897
rect 128529 281835 128839 281869
rect 128529 281807 128577 281835
rect 128605 281807 128639 281835
rect 128667 281807 128701 281835
rect 128729 281807 128763 281835
rect 128791 281807 128839 281835
rect 128529 281773 128839 281807
rect 128529 281745 128577 281773
rect 128605 281745 128639 281773
rect 128667 281745 128701 281773
rect 128729 281745 128763 281773
rect 128791 281745 128839 281773
rect 128529 272959 128839 281745
rect 128529 272931 128577 272959
rect 128605 272931 128639 272959
rect 128667 272931 128701 272959
rect 128729 272931 128763 272959
rect 128791 272931 128839 272959
rect 128529 272897 128839 272931
rect 128529 272869 128577 272897
rect 128605 272869 128639 272897
rect 128667 272869 128701 272897
rect 128729 272869 128763 272897
rect 128791 272869 128839 272897
rect 128529 272835 128839 272869
rect 128529 272807 128577 272835
rect 128605 272807 128639 272835
rect 128667 272807 128701 272835
rect 128729 272807 128763 272835
rect 128791 272807 128839 272835
rect 128529 272773 128839 272807
rect 128529 272745 128577 272773
rect 128605 272745 128639 272773
rect 128667 272745 128701 272773
rect 128729 272745 128763 272773
rect 128791 272745 128839 272773
rect 128529 263959 128839 272745
rect 128529 263931 128577 263959
rect 128605 263931 128639 263959
rect 128667 263931 128701 263959
rect 128729 263931 128763 263959
rect 128791 263931 128839 263959
rect 128529 263897 128839 263931
rect 128529 263869 128577 263897
rect 128605 263869 128639 263897
rect 128667 263869 128701 263897
rect 128729 263869 128763 263897
rect 128791 263869 128839 263897
rect 128529 263835 128839 263869
rect 128529 263807 128577 263835
rect 128605 263807 128639 263835
rect 128667 263807 128701 263835
rect 128729 263807 128763 263835
rect 128791 263807 128839 263835
rect 128529 263773 128839 263807
rect 128529 263745 128577 263773
rect 128605 263745 128639 263773
rect 128667 263745 128701 263773
rect 128729 263745 128763 263773
rect 128791 263745 128839 263773
rect 128529 254959 128839 263745
rect 128529 254931 128577 254959
rect 128605 254931 128639 254959
rect 128667 254931 128701 254959
rect 128729 254931 128763 254959
rect 128791 254931 128839 254959
rect 128529 254897 128839 254931
rect 128529 254869 128577 254897
rect 128605 254869 128639 254897
rect 128667 254869 128701 254897
rect 128729 254869 128763 254897
rect 128791 254869 128839 254897
rect 128529 254835 128839 254869
rect 128529 254807 128577 254835
rect 128605 254807 128639 254835
rect 128667 254807 128701 254835
rect 128729 254807 128763 254835
rect 128791 254807 128839 254835
rect 128529 254773 128839 254807
rect 128529 254745 128577 254773
rect 128605 254745 128639 254773
rect 128667 254745 128701 254773
rect 128729 254745 128763 254773
rect 128791 254745 128839 254773
rect 128529 254075 128839 254745
rect 130389 299670 130699 299718
rect 130389 299642 130437 299670
rect 130465 299642 130499 299670
rect 130527 299642 130561 299670
rect 130589 299642 130623 299670
rect 130651 299642 130699 299670
rect 130389 299608 130699 299642
rect 130389 299580 130437 299608
rect 130465 299580 130499 299608
rect 130527 299580 130561 299608
rect 130589 299580 130623 299608
rect 130651 299580 130699 299608
rect 130389 299546 130699 299580
rect 130389 299518 130437 299546
rect 130465 299518 130499 299546
rect 130527 299518 130561 299546
rect 130589 299518 130623 299546
rect 130651 299518 130699 299546
rect 130389 299484 130699 299518
rect 130389 299456 130437 299484
rect 130465 299456 130499 299484
rect 130527 299456 130561 299484
rect 130589 299456 130623 299484
rect 130651 299456 130699 299484
rect 130389 293959 130699 299456
rect 130389 293931 130437 293959
rect 130465 293931 130499 293959
rect 130527 293931 130561 293959
rect 130589 293931 130623 293959
rect 130651 293931 130699 293959
rect 130389 293897 130699 293931
rect 130389 293869 130437 293897
rect 130465 293869 130499 293897
rect 130527 293869 130561 293897
rect 130589 293869 130623 293897
rect 130651 293869 130699 293897
rect 130389 293835 130699 293869
rect 130389 293807 130437 293835
rect 130465 293807 130499 293835
rect 130527 293807 130561 293835
rect 130589 293807 130623 293835
rect 130651 293807 130699 293835
rect 130389 293773 130699 293807
rect 130389 293745 130437 293773
rect 130465 293745 130499 293773
rect 130527 293745 130561 293773
rect 130589 293745 130623 293773
rect 130651 293745 130699 293773
rect 130389 284959 130699 293745
rect 130389 284931 130437 284959
rect 130465 284931 130499 284959
rect 130527 284931 130561 284959
rect 130589 284931 130623 284959
rect 130651 284931 130699 284959
rect 130389 284897 130699 284931
rect 130389 284869 130437 284897
rect 130465 284869 130499 284897
rect 130527 284869 130561 284897
rect 130589 284869 130623 284897
rect 130651 284869 130699 284897
rect 130389 284835 130699 284869
rect 130389 284807 130437 284835
rect 130465 284807 130499 284835
rect 130527 284807 130561 284835
rect 130589 284807 130623 284835
rect 130651 284807 130699 284835
rect 130389 284773 130699 284807
rect 130389 284745 130437 284773
rect 130465 284745 130499 284773
rect 130527 284745 130561 284773
rect 130589 284745 130623 284773
rect 130651 284745 130699 284773
rect 130389 275959 130699 284745
rect 130389 275931 130437 275959
rect 130465 275931 130499 275959
rect 130527 275931 130561 275959
rect 130589 275931 130623 275959
rect 130651 275931 130699 275959
rect 130389 275897 130699 275931
rect 130389 275869 130437 275897
rect 130465 275869 130499 275897
rect 130527 275869 130561 275897
rect 130589 275869 130623 275897
rect 130651 275869 130699 275897
rect 130389 275835 130699 275869
rect 130389 275807 130437 275835
rect 130465 275807 130499 275835
rect 130527 275807 130561 275835
rect 130589 275807 130623 275835
rect 130651 275807 130699 275835
rect 130389 275773 130699 275807
rect 130389 275745 130437 275773
rect 130465 275745 130499 275773
rect 130527 275745 130561 275773
rect 130589 275745 130623 275773
rect 130651 275745 130699 275773
rect 130389 266959 130699 275745
rect 130389 266931 130437 266959
rect 130465 266931 130499 266959
rect 130527 266931 130561 266959
rect 130589 266931 130623 266959
rect 130651 266931 130699 266959
rect 130389 266897 130699 266931
rect 130389 266869 130437 266897
rect 130465 266869 130499 266897
rect 130527 266869 130561 266897
rect 130589 266869 130623 266897
rect 130651 266869 130699 266897
rect 130389 266835 130699 266869
rect 130389 266807 130437 266835
rect 130465 266807 130499 266835
rect 130527 266807 130561 266835
rect 130589 266807 130623 266835
rect 130651 266807 130699 266835
rect 130389 266773 130699 266807
rect 130389 266745 130437 266773
rect 130465 266745 130499 266773
rect 130527 266745 130561 266773
rect 130589 266745 130623 266773
rect 130651 266745 130699 266773
rect 130389 257959 130699 266745
rect 130389 257931 130437 257959
rect 130465 257931 130499 257959
rect 130527 257931 130561 257959
rect 130589 257931 130623 257959
rect 130651 257931 130699 257959
rect 130389 257897 130699 257931
rect 130389 257869 130437 257897
rect 130465 257869 130499 257897
rect 130527 257869 130561 257897
rect 130589 257869 130623 257897
rect 130651 257869 130699 257897
rect 130389 257835 130699 257869
rect 130389 257807 130437 257835
rect 130465 257807 130499 257835
rect 130527 257807 130561 257835
rect 130589 257807 130623 257835
rect 130651 257807 130699 257835
rect 130389 257773 130699 257807
rect 130389 257745 130437 257773
rect 130465 257745 130499 257773
rect 130527 257745 130561 257773
rect 130589 257745 130623 257773
rect 130651 257745 130699 257773
rect 130389 254075 130699 257745
rect 137529 299190 137839 299718
rect 137529 299162 137577 299190
rect 137605 299162 137639 299190
rect 137667 299162 137701 299190
rect 137729 299162 137763 299190
rect 137791 299162 137839 299190
rect 137529 299128 137839 299162
rect 137529 299100 137577 299128
rect 137605 299100 137639 299128
rect 137667 299100 137701 299128
rect 137729 299100 137763 299128
rect 137791 299100 137839 299128
rect 137529 299066 137839 299100
rect 137529 299038 137577 299066
rect 137605 299038 137639 299066
rect 137667 299038 137701 299066
rect 137729 299038 137763 299066
rect 137791 299038 137839 299066
rect 137529 299004 137839 299038
rect 137529 298976 137577 299004
rect 137605 298976 137639 299004
rect 137667 298976 137701 299004
rect 137729 298976 137763 299004
rect 137791 298976 137839 299004
rect 137529 290959 137839 298976
rect 137529 290931 137577 290959
rect 137605 290931 137639 290959
rect 137667 290931 137701 290959
rect 137729 290931 137763 290959
rect 137791 290931 137839 290959
rect 137529 290897 137839 290931
rect 137529 290869 137577 290897
rect 137605 290869 137639 290897
rect 137667 290869 137701 290897
rect 137729 290869 137763 290897
rect 137791 290869 137839 290897
rect 137529 290835 137839 290869
rect 137529 290807 137577 290835
rect 137605 290807 137639 290835
rect 137667 290807 137701 290835
rect 137729 290807 137763 290835
rect 137791 290807 137839 290835
rect 137529 290773 137839 290807
rect 137529 290745 137577 290773
rect 137605 290745 137639 290773
rect 137667 290745 137701 290773
rect 137729 290745 137763 290773
rect 137791 290745 137839 290773
rect 137529 281959 137839 290745
rect 137529 281931 137577 281959
rect 137605 281931 137639 281959
rect 137667 281931 137701 281959
rect 137729 281931 137763 281959
rect 137791 281931 137839 281959
rect 137529 281897 137839 281931
rect 137529 281869 137577 281897
rect 137605 281869 137639 281897
rect 137667 281869 137701 281897
rect 137729 281869 137763 281897
rect 137791 281869 137839 281897
rect 137529 281835 137839 281869
rect 137529 281807 137577 281835
rect 137605 281807 137639 281835
rect 137667 281807 137701 281835
rect 137729 281807 137763 281835
rect 137791 281807 137839 281835
rect 137529 281773 137839 281807
rect 137529 281745 137577 281773
rect 137605 281745 137639 281773
rect 137667 281745 137701 281773
rect 137729 281745 137763 281773
rect 137791 281745 137839 281773
rect 137529 272959 137839 281745
rect 137529 272931 137577 272959
rect 137605 272931 137639 272959
rect 137667 272931 137701 272959
rect 137729 272931 137763 272959
rect 137791 272931 137839 272959
rect 137529 272897 137839 272931
rect 137529 272869 137577 272897
rect 137605 272869 137639 272897
rect 137667 272869 137701 272897
rect 137729 272869 137763 272897
rect 137791 272869 137839 272897
rect 137529 272835 137839 272869
rect 137529 272807 137577 272835
rect 137605 272807 137639 272835
rect 137667 272807 137701 272835
rect 137729 272807 137763 272835
rect 137791 272807 137839 272835
rect 137529 272773 137839 272807
rect 137529 272745 137577 272773
rect 137605 272745 137639 272773
rect 137667 272745 137701 272773
rect 137729 272745 137763 272773
rect 137791 272745 137839 272773
rect 137529 263959 137839 272745
rect 137529 263931 137577 263959
rect 137605 263931 137639 263959
rect 137667 263931 137701 263959
rect 137729 263931 137763 263959
rect 137791 263931 137839 263959
rect 137529 263897 137839 263931
rect 137529 263869 137577 263897
rect 137605 263869 137639 263897
rect 137667 263869 137701 263897
rect 137729 263869 137763 263897
rect 137791 263869 137839 263897
rect 137529 263835 137839 263869
rect 137529 263807 137577 263835
rect 137605 263807 137639 263835
rect 137667 263807 137701 263835
rect 137729 263807 137763 263835
rect 137791 263807 137839 263835
rect 137529 263773 137839 263807
rect 137529 263745 137577 263773
rect 137605 263745 137639 263773
rect 137667 263745 137701 263773
rect 137729 263745 137763 263773
rect 137791 263745 137839 263773
rect 137529 254959 137839 263745
rect 137529 254931 137577 254959
rect 137605 254931 137639 254959
rect 137667 254931 137701 254959
rect 137729 254931 137763 254959
rect 137791 254931 137839 254959
rect 137529 254897 137839 254931
rect 137529 254869 137577 254897
rect 137605 254869 137639 254897
rect 137667 254869 137701 254897
rect 137729 254869 137763 254897
rect 137791 254869 137839 254897
rect 137529 254835 137839 254869
rect 137529 254807 137577 254835
rect 137605 254807 137639 254835
rect 137667 254807 137701 254835
rect 137729 254807 137763 254835
rect 137791 254807 137839 254835
rect 137529 254773 137839 254807
rect 137529 254745 137577 254773
rect 137605 254745 137639 254773
rect 137667 254745 137701 254773
rect 137729 254745 137763 254773
rect 137791 254745 137839 254773
rect 137529 254075 137839 254745
rect 139389 299670 139699 299718
rect 139389 299642 139437 299670
rect 139465 299642 139499 299670
rect 139527 299642 139561 299670
rect 139589 299642 139623 299670
rect 139651 299642 139699 299670
rect 139389 299608 139699 299642
rect 139389 299580 139437 299608
rect 139465 299580 139499 299608
rect 139527 299580 139561 299608
rect 139589 299580 139623 299608
rect 139651 299580 139699 299608
rect 139389 299546 139699 299580
rect 139389 299518 139437 299546
rect 139465 299518 139499 299546
rect 139527 299518 139561 299546
rect 139589 299518 139623 299546
rect 139651 299518 139699 299546
rect 139389 299484 139699 299518
rect 139389 299456 139437 299484
rect 139465 299456 139499 299484
rect 139527 299456 139561 299484
rect 139589 299456 139623 299484
rect 139651 299456 139699 299484
rect 139389 293959 139699 299456
rect 139389 293931 139437 293959
rect 139465 293931 139499 293959
rect 139527 293931 139561 293959
rect 139589 293931 139623 293959
rect 139651 293931 139699 293959
rect 139389 293897 139699 293931
rect 139389 293869 139437 293897
rect 139465 293869 139499 293897
rect 139527 293869 139561 293897
rect 139589 293869 139623 293897
rect 139651 293869 139699 293897
rect 139389 293835 139699 293869
rect 139389 293807 139437 293835
rect 139465 293807 139499 293835
rect 139527 293807 139561 293835
rect 139589 293807 139623 293835
rect 139651 293807 139699 293835
rect 139389 293773 139699 293807
rect 139389 293745 139437 293773
rect 139465 293745 139499 293773
rect 139527 293745 139561 293773
rect 139589 293745 139623 293773
rect 139651 293745 139699 293773
rect 139389 284959 139699 293745
rect 139389 284931 139437 284959
rect 139465 284931 139499 284959
rect 139527 284931 139561 284959
rect 139589 284931 139623 284959
rect 139651 284931 139699 284959
rect 139389 284897 139699 284931
rect 139389 284869 139437 284897
rect 139465 284869 139499 284897
rect 139527 284869 139561 284897
rect 139589 284869 139623 284897
rect 139651 284869 139699 284897
rect 139389 284835 139699 284869
rect 139389 284807 139437 284835
rect 139465 284807 139499 284835
rect 139527 284807 139561 284835
rect 139589 284807 139623 284835
rect 139651 284807 139699 284835
rect 139389 284773 139699 284807
rect 139389 284745 139437 284773
rect 139465 284745 139499 284773
rect 139527 284745 139561 284773
rect 139589 284745 139623 284773
rect 139651 284745 139699 284773
rect 139389 275959 139699 284745
rect 139389 275931 139437 275959
rect 139465 275931 139499 275959
rect 139527 275931 139561 275959
rect 139589 275931 139623 275959
rect 139651 275931 139699 275959
rect 139389 275897 139699 275931
rect 139389 275869 139437 275897
rect 139465 275869 139499 275897
rect 139527 275869 139561 275897
rect 139589 275869 139623 275897
rect 139651 275869 139699 275897
rect 139389 275835 139699 275869
rect 139389 275807 139437 275835
rect 139465 275807 139499 275835
rect 139527 275807 139561 275835
rect 139589 275807 139623 275835
rect 139651 275807 139699 275835
rect 139389 275773 139699 275807
rect 139389 275745 139437 275773
rect 139465 275745 139499 275773
rect 139527 275745 139561 275773
rect 139589 275745 139623 275773
rect 139651 275745 139699 275773
rect 139389 266959 139699 275745
rect 139389 266931 139437 266959
rect 139465 266931 139499 266959
rect 139527 266931 139561 266959
rect 139589 266931 139623 266959
rect 139651 266931 139699 266959
rect 139389 266897 139699 266931
rect 139389 266869 139437 266897
rect 139465 266869 139499 266897
rect 139527 266869 139561 266897
rect 139589 266869 139623 266897
rect 139651 266869 139699 266897
rect 139389 266835 139699 266869
rect 139389 266807 139437 266835
rect 139465 266807 139499 266835
rect 139527 266807 139561 266835
rect 139589 266807 139623 266835
rect 139651 266807 139699 266835
rect 139389 266773 139699 266807
rect 139389 266745 139437 266773
rect 139465 266745 139499 266773
rect 139527 266745 139561 266773
rect 139589 266745 139623 266773
rect 139651 266745 139699 266773
rect 139389 257959 139699 266745
rect 139389 257931 139437 257959
rect 139465 257931 139499 257959
rect 139527 257931 139561 257959
rect 139589 257931 139623 257959
rect 139651 257931 139699 257959
rect 139389 257897 139699 257931
rect 139389 257869 139437 257897
rect 139465 257869 139499 257897
rect 139527 257869 139561 257897
rect 139589 257869 139623 257897
rect 139651 257869 139699 257897
rect 139389 257835 139699 257869
rect 139389 257807 139437 257835
rect 139465 257807 139499 257835
rect 139527 257807 139561 257835
rect 139589 257807 139623 257835
rect 139651 257807 139699 257835
rect 139389 257773 139699 257807
rect 139389 257745 139437 257773
rect 139465 257745 139499 257773
rect 139527 257745 139561 257773
rect 139589 257745 139623 257773
rect 139651 257745 139699 257773
rect 139389 254075 139699 257745
rect 146529 299190 146839 299718
rect 146529 299162 146577 299190
rect 146605 299162 146639 299190
rect 146667 299162 146701 299190
rect 146729 299162 146763 299190
rect 146791 299162 146839 299190
rect 146529 299128 146839 299162
rect 146529 299100 146577 299128
rect 146605 299100 146639 299128
rect 146667 299100 146701 299128
rect 146729 299100 146763 299128
rect 146791 299100 146839 299128
rect 146529 299066 146839 299100
rect 146529 299038 146577 299066
rect 146605 299038 146639 299066
rect 146667 299038 146701 299066
rect 146729 299038 146763 299066
rect 146791 299038 146839 299066
rect 146529 299004 146839 299038
rect 146529 298976 146577 299004
rect 146605 298976 146639 299004
rect 146667 298976 146701 299004
rect 146729 298976 146763 299004
rect 146791 298976 146839 299004
rect 146529 290959 146839 298976
rect 146529 290931 146577 290959
rect 146605 290931 146639 290959
rect 146667 290931 146701 290959
rect 146729 290931 146763 290959
rect 146791 290931 146839 290959
rect 146529 290897 146839 290931
rect 146529 290869 146577 290897
rect 146605 290869 146639 290897
rect 146667 290869 146701 290897
rect 146729 290869 146763 290897
rect 146791 290869 146839 290897
rect 146529 290835 146839 290869
rect 146529 290807 146577 290835
rect 146605 290807 146639 290835
rect 146667 290807 146701 290835
rect 146729 290807 146763 290835
rect 146791 290807 146839 290835
rect 146529 290773 146839 290807
rect 146529 290745 146577 290773
rect 146605 290745 146639 290773
rect 146667 290745 146701 290773
rect 146729 290745 146763 290773
rect 146791 290745 146839 290773
rect 146529 281959 146839 290745
rect 146529 281931 146577 281959
rect 146605 281931 146639 281959
rect 146667 281931 146701 281959
rect 146729 281931 146763 281959
rect 146791 281931 146839 281959
rect 146529 281897 146839 281931
rect 146529 281869 146577 281897
rect 146605 281869 146639 281897
rect 146667 281869 146701 281897
rect 146729 281869 146763 281897
rect 146791 281869 146839 281897
rect 146529 281835 146839 281869
rect 146529 281807 146577 281835
rect 146605 281807 146639 281835
rect 146667 281807 146701 281835
rect 146729 281807 146763 281835
rect 146791 281807 146839 281835
rect 146529 281773 146839 281807
rect 146529 281745 146577 281773
rect 146605 281745 146639 281773
rect 146667 281745 146701 281773
rect 146729 281745 146763 281773
rect 146791 281745 146839 281773
rect 146529 272959 146839 281745
rect 146529 272931 146577 272959
rect 146605 272931 146639 272959
rect 146667 272931 146701 272959
rect 146729 272931 146763 272959
rect 146791 272931 146839 272959
rect 146529 272897 146839 272931
rect 146529 272869 146577 272897
rect 146605 272869 146639 272897
rect 146667 272869 146701 272897
rect 146729 272869 146763 272897
rect 146791 272869 146839 272897
rect 146529 272835 146839 272869
rect 146529 272807 146577 272835
rect 146605 272807 146639 272835
rect 146667 272807 146701 272835
rect 146729 272807 146763 272835
rect 146791 272807 146839 272835
rect 146529 272773 146839 272807
rect 146529 272745 146577 272773
rect 146605 272745 146639 272773
rect 146667 272745 146701 272773
rect 146729 272745 146763 272773
rect 146791 272745 146839 272773
rect 146529 263959 146839 272745
rect 146529 263931 146577 263959
rect 146605 263931 146639 263959
rect 146667 263931 146701 263959
rect 146729 263931 146763 263959
rect 146791 263931 146839 263959
rect 146529 263897 146839 263931
rect 146529 263869 146577 263897
rect 146605 263869 146639 263897
rect 146667 263869 146701 263897
rect 146729 263869 146763 263897
rect 146791 263869 146839 263897
rect 146529 263835 146839 263869
rect 146529 263807 146577 263835
rect 146605 263807 146639 263835
rect 146667 263807 146701 263835
rect 146729 263807 146763 263835
rect 146791 263807 146839 263835
rect 146529 263773 146839 263807
rect 146529 263745 146577 263773
rect 146605 263745 146639 263773
rect 146667 263745 146701 263773
rect 146729 263745 146763 263773
rect 146791 263745 146839 263773
rect 146529 254959 146839 263745
rect 146529 254931 146577 254959
rect 146605 254931 146639 254959
rect 146667 254931 146701 254959
rect 146729 254931 146763 254959
rect 146791 254931 146839 254959
rect 146529 254897 146839 254931
rect 146529 254869 146577 254897
rect 146605 254869 146639 254897
rect 146667 254869 146701 254897
rect 146729 254869 146763 254897
rect 146791 254869 146839 254897
rect 146529 254835 146839 254869
rect 146529 254807 146577 254835
rect 146605 254807 146639 254835
rect 146667 254807 146701 254835
rect 146729 254807 146763 254835
rect 146791 254807 146839 254835
rect 146529 254773 146839 254807
rect 146529 254745 146577 254773
rect 146605 254745 146639 254773
rect 146667 254745 146701 254773
rect 146729 254745 146763 254773
rect 146791 254745 146839 254773
rect 146529 254075 146839 254745
rect 148389 299670 148699 299718
rect 148389 299642 148437 299670
rect 148465 299642 148499 299670
rect 148527 299642 148561 299670
rect 148589 299642 148623 299670
rect 148651 299642 148699 299670
rect 148389 299608 148699 299642
rect 148389 299580 148437 299608
rect 148465 299580 148499 299608
rect 148527 299580 148561 299608
rect 148589 299580 148623 299608
rect 148651 299580 148699 299608
rect 148389 299546 148699 299580
rect 148389 299518 148437 299546
rect 148465 299518 148499 299546
rect 148527 299518 148561 299546
rect 148589 299518 148623 299546
rect 148651 299518 148699 299546
rect 148389 299484 148699 299518
rect 148389 299456 148437 299484
rect 148465 299456 148499 299484
rect 148527 299456 148561 299484
rect 148589 299456 148623 299484
rect 148651 299456 148699 299484
rect 148389 293959 148699 299456
rect 148389 293931 148437 293959
rect 148465 293931 148499 293959
rect 148527 293931 148561 293959
rect 148589 293931 148623 293959
rect 148651 293931 148699 293959
rect 148389 293897 148699 293931
rect 148389 293869 148437 293897
rect 148465 293869 148499 293897
rect 148527 293869 148561 293897
rect 148589 293869 148623 293897
rect 148651 293869 148699 293897
rect 148389 293835 148699 293869
rect 148389 293807 148437 293835
rect 148465 293807 148499 293835
rect 148527 293807 148561 293835
rect 148589 293807 148623 293835
rect 148651 293807 148699 293835
rect 148389 293773 148699 293807
rect 148389 293745 148437 293773
rect 148465 293745 148499 293773
rect 148527 293745 148561 293773
rect 148589 293745 148623 293773
rect 148651 293745 148699 293773
rect 148389 284959 148699 293745
rect 148389 284931 148437 284959
rect 148465 284931 148499 284959
rect 148527 284931 148561 284959
rect 148589 284931 148623 284959
rect 148651 284931 148699 284959
rect 148389 284897 148699 284931
rect 148389 284869 148437 284897
rect 148465 284869 148499 284897
rect 148527 284869 148561 284897
rect 148589 284869 148623 284897
rect 148651 284869 148699 284897
rect 148389 284835 148699 284869
rect 148389 284807 148437 284835
rect 148465 284807 148499 284835
rect 148527 284807 148561 284835
rect 148589 284807 148623 284835
rect 148651 284807 148699 284835
rect 148389 284773 148699 284807
rect 148389 284745 148437 284773
rect 148465 284745 148499 284773
rect 148527 284745 148561 284773
rect 148589 284745 148623 284773
rect 148651 284745 148699 284773
rect 148389 275959 148699 284745
rect 148389 275931 148437 275959
rect 148465 275931 148499 275959
rect 148527 275931 148561 275959
rect 148589 275931 148623 275959
rect 148651 275931 148699 275959
rect 148389 275897 148699 275931
rect 148389 275869 148437 275897
rect 148465 275869 148499 275897
rect 148527 275869 148561 275897
rect 148589 275869 148623 275897
rect 148651 275869 148699 275897
rect 148389 275835 148699 275869
rect 148389 275807 148437 275835
rect 148465 275807 148499 275835
rect 148527 275807 148561 275835
rect 148589 275807 148623 275835
rect 148651 275807 148699 275835
rect 148389 275773 148699 275807
rect 148389 275745 148437 275773
rect 148465 275745 148499 275773
rect 148527 275745 148561 275773
rect 148589 275745 148623 275773
rect 148651 275745 148699 275773
rect 148389 266959 148699 275745
rect 148389 266931 148437 266959
rect 148465 266931 148499 266959
rect 148527 266931 148561 266959
rect 148589 266931 148623 266959
rect 148651 266931 148699 266959
rect 148389 266897 148699 266931
rect 148389 266869 148437 266897
rect 148465 266869 148499 266897
rect 148527 266869 148561 266897
rect 148589 266869 148623 266897
rect 148651 266869 148699 266897
rect 148389 266835 148699 266869
rect 148389 266807 148437 266835
rect 148465 266807 148499 266835
rect 148527 266807 148561 266835
rect 148589 266807 148623 266835
rect 148651 266807 148699 266835
rect 148389 266773 148699 266807
rect 148389 266745 148437 266773
rect 148465 266745 148499 266773
rect 148527 266745 148561 266773
rect 148589 266745 148623 266773
rect 148651 266745 148699 266773
rect 148389 257959 148699 266745
rect 148389 257931 148437 257959
rect 148465 257931 148499 257959
rect 148527 257931 148561 257959
rect 148589 257931 148623 257959
rect 148651 257931 148699 257959
rect 148389 257897 148699 257931
rect 148389 257869 148437 257897
rect 148465 257869 148499 257897
rect 148527 257869 148561 257897
rect 148589 257869 148623 257897
rect 148651 257869 148699 257897
rect 148389 257835 148699 257869
rect 148389 257807 148437 257835
rect 148465 257807 148499 257835
rect 148527 257807 148561 257835
rect 148589 257807 148623 257835
rect 148651 257807 148699 257835
rect 148389 257773 148699 257807
rect 148389 257745 148437 257773
rect 148465 257745 148499 257773
rect 148527 257745 148561 257773
rect 148589 257745 148623 257773
rect 148651 257745 148699 257773
rect 148389 254075 148699 257745
rect 155529 299190 155839 299718
rect 155529 299162 155577 299190
rect 155605 299162 155639 299190
rect 155667 299162 155701 299190
rect 155729 299162 155763 299190
rect 155791 299162 155839 299190
rect 155529 299128 155839 299162
rect 155529 299100 155577 299128
rect 155605 299100 155639 299128
rect 155667 299100 155701 299128
rect 155729 299100 155763 299128
rect 155791 299100 155839 299128
rect 155529 299066 155839 299100
rect 155529 299038 155577 299066
rect 155605 299038 155639 299066
rect 155667 299038 155701 299066
rect 155729 299038 155763 299066
rect 155791 299038 155839 299066
rect 155529 299004 155839 299038
rect 155529 298976 155577 299004
rect 155605 298976 155639 299004
rect 155667 298976 155701 299004
rect 155729 298976 155763 299004
rect 155791 298976 155839 299004
rect 155529 290959 155839 298976
rect 155529 290931 155577 290959
rect 155605 290931 155639 290959
rect 155667 290931 155701 290959
rect 155729 290931 155763 290959
rect 155791 290931 155839 290959
rect 155529 290897 155839 290931
rect 155529 290869 155577 290897
rect 155605 290869 155639 290897
rect 155667 290869 155701 290897
rect 155729 290869 155763 290897
rect 155791 290869 155839 290897
rect 155529 290835 155839 290869
rect 155529 290807 155577 290835
rect 155605 290807 155639 290835
rect 155667 290807 155701 290835
rect 155729 290807 155763 290835
rect 155791 290807 155839 290835
rect 155529 290773 155839 290807
rect 155529 290745 155577 290773
rect 155605 290745 155639 290773
rect 155667 290745 155701 290773
rect 155729 290745 155763 290773
rect 155791 290745 155839 290773
rect 155529 281959 155839 290745
rect 155529 281931 155577 281959
rect 155605 281931 155639 281959
rect 155667 281931 155701 281959
rect 155729 281931 155763 281959
rect 155791 281931 155839 281959
rect 155529 281897 155839 281931
rect 155529 281869 155577 281897
rect 155605 281869 155639 281897
rect 155667 281869 155701 281897
rect 155729 281869 155763 281897
rect 155791 281869 155839 281897
rect 155529 281835 155839 281869
rect 155529 281807 155577 281835
rect 155605 281807 155639 281835
rect 155667 281807 155701 281835
rect 155729 281807 155763 281835
rect 155791 281807 155839 281835
rect 155529 281773 155839 281807
rect 155529 281745 155577 281773
rect 155605 281745 155639 281773
rect 155667 281745 155701 281773
rect 155729 281745 155763 281773
rect 155791 281745 155839 281773
rect 155529 272959 155839 281745
rect 155529 272931 155577 272959
rect 155605 272931 155639 272959
rect 155667 272931 155701 272959
rect 155729 272931 155763 272959
rect 155791 272931 155839 272959
rect 155529 272897 155839 272931
rect 155529 272869 155577 272897
rect 155605 272869 155639 272897
rect 155667 272869 155701 272897
rect 155729 272869 155763 272897
rect 155791 272869 155839 272897
rect 155529 272835 155839 272869
rect 155529 272807 155577 272835
rect 155605 272807 155639 272835
rect 155667 272807 155701 272835
rect 155729 272807 155763 272835
rect 155791 272807 155839 272835
rect 155529 272773 155839 272807
rect 155529 272745 155577 272773
rect 155605 272745 155639 272773
rect 155667 272745 155701 272773
rect 155729 272745 155763 272773
rect 155791 272745 155839 272773
rect 155529 263959 155839 272745
rect 155529 263931 155577 263959
rect 155605 263931 155639 263959
rect 155667 263931 155701 263959
rect 155729 263931 155763 263959
rect 155791 263931 155839 263959
rect 155529 263897 155839 263931
rect 155529 263869 155577 263897
rect 155605 263869 155639 263897
rect 155667 263869 155701 263897
rect 155729 263869 155763 263897
rect 155791 263869 155839 263897
rect 155529 263835 155839 263869
rect 155529 263807 155577 263835
rect 155605 263807 155639 263835
rect 155667 263807 155701 263835
rect 155729 263807 155763 263835
rect 155791 263807 155839 263835
rect 155529 263773 155839 263807
rect 155529 263745 155577 263773
rect 155605 263745 155639 263773
rect 155667 263745 155701 263773
rect 155729 263745 155763 263773
rect 155791 263745 155839 263773
rect 155529 254959 155839 263745
rect 155529 254931 155577 254959
rect 155605 254931 155639 254959
rect 155667 254931 155701 254959
rect 155729 254931 155763 254959
rect 155791 254931 155839 254959
rect 155529 254897 155839 254931
rect 155529 254869 155577 254897
rect 155605 254869 155639 254897
rect 155667 254869 155701 254897
rect 155729 254869 155763 254897
rect 155791 254869 155839 254897
rect 155529 254835 155839 254869
rect 155529 254807 155577 254835
rect 155605 254807 155639 254835
rect 155667 254807 155701 254835
rect 155729 254807 155763 254835
rect 155791 254807 155839 254835
rect 155529 254773 155839 254807
rect 155529 254745 155577 254773
rect 155605 254745 155639 254773
rect 155667 254745 155701 254773
rect 155729 254745 155763 254773
rect 155791 254745 155839 254773
rect 155529 254394 155839 254745
rect 157389 299670 157699 299718
rect 157389 299642 157437 299670
rect 157465 299642 157499 299670
rect 157527 299642 157561 299670
rect 157589 299642 157623 299670
rect 157651 299642 157699 299670
rect 157389 299608 157699 299642
rect 157389 299580 157437 299608
rect 157465 299580 157499 299608
rect 157527 299580 157561 299608
rect 157589 299580 157623 299608
rect 157651 299580 157699 299608
rect 157389 299546 157699 299580
rect 157389 299518 157437 299546
rect 157465 299518 157499 299546
rect 157527 299518 157561 299546
rect 157589 299518 157623 299546
rect 157651 299518 157699 299546
rect 157389 299484 157699 299518
rect 157389 299456 157437 299484
rect 157465 299456 157499 299484
rect 157527 299456 157561 299484
rect 157589 299456 157623 299484
rect 157651 299456 157699 299484
rect 157389 293959 157699 299456
rect 157389 293931 157437 293959
rect 157465 293931 157499 293959
rect 157527 293931 157561 293959
rect 157589 293931 157623 293959
rect 157651 293931 157699 293959
rect 157389 293897 157699 293931
rect 157389 293869 157437 293897
rect 157465 293869 157499 293897
rect 157527 293869 157561 293897
rect 157589 293869 157623 293897
rect 157651 293869 157699 293897
rect 157389 293835 157699 293869
rect 157389 293807 157437 293835
rect 157465 293807 157499 293835
rect 157527 293807 157561 293835
rect 157589 293807 157623 293835
rect 157651 293807 157699 293835
rect 157389 293773 157699 293807
rect 157389 293745 157437 293773
rect 157465 293745 157499 293773
rect 157527 293745 157561 293773
rect 157589 293745 157623 293773
rect 157651 293745 157699 293773
rect 157389 284959 157699 293745
rect 157389 284931 157437 284959
rect 157465 284931 157499 284959
rect 157527 284931 157561 284959
rect 157589 284931 157623 284959
rect 157651 284931 157699 284959
rect 157389 284897 157699 284931
rect 157389 284869 157437 284897
rect 157465 284869 157499 284897
rect 157527 284869 157561 284897
rect 157589 284869 157623 284897
rect 157651 284869 157699 284897
rect 157389 284835 157699 284869
rect 157389 284807 157437 284835
rect 157465 284807 157499 284835
rect 157527 284807 157561 284835
rect 157589 284807 157623 284835
rect 157651 284807 157699 284835
rect 157389 284773 157699 284807
rect 157389 284745 157437 284773
rect 157465 284745 157499 284773
rect 157527 284745 157561 284773
rect 157589 284745 157623 284773
rect 157651 284745 157699 284773
rect 157389 275959 157699 284745
rect 157389 275931 157437 275959
rect 157465 275931 157499 275959
rect 157527 275931 157561 275959
rect 157589 275931 157623 275959
rect 157651 275931 157699 275959
rect 157389 275897 157699 275931
rect 157389 275869 157437 275897
rect 157465 275869 157499 275897
rect 157527 275869 157561 275897
rect 157589 275869 157623 275897
rect 157651 275869 157699 275897
rect 157389 275835 157699 275869
rect 157389 275807 157437 275835
rect 157465 275807 157499 275835
rect 157527 275807 157561 275835
rect 157589 275807 157623 275835
rect 157651 275807 157699 275835
rect 157389 275773 157699 275807
rect 157389 275745 157437 275773
rect 157465 275745 157499 275773
rect 157527 275745 157561 275773
rect 157589 275745 157623 275773
rect 157651 275745 157699 275773
rect 157389 266959 157699 275745
rect 157389 266931 157437 266959
rect 157465 266931 157499 266959
rect 157527 266931 157561 266959
rect 157589 266931 157623 266959
rect 157651 266931 157699 266959
rect 157389 266897 157699 266931
rect 157389 266869 157437 266897
rect 157465 266869 157499 266897
rect 157527 266869 157561 266897
rect 157589 266869 157623 266897
rect 157651 266869 157699 266897
rect 157389 266835 157699 266869
rect 157389 266807 157437 266835
rect 157465 266807 157499 266835
rect 157527 266807 157561 266835
rect 157589 266807 157623 266835
rect 157651 266807 157699 266835
rect 157389 266773 157699 266807
rect 157389 266745 157437 266773
rect 157465 266745 157499 266773
rect 157527 266745 157561 266773
rect 157589 266745 157623 266773
rect 157651 266745 157699 266773
rect 157389 257959 157699 266745
rect 157389 257931 157437 257959
rect 157465 257931 157499 257959
rect 157527 257931 157561 257959
rect 157589 257931 157623 257959
rect 157651 257931 157699 257959
rect 157389 257897 157699 257931
rect 157389 257869 157437 257897
rect 157465 257869 157499 257897
rect 157527 257869 157561 257897
rect 157589 257869 157623 257897
rect 157651 257869 157699 257897
rect 157389 257835 157699 257869
rect 157389 257807 157437 257835
rect 157465 257807 157499 257835
rect 157527 257807 157561 257835
rect 157589 257807 157623 257835
rect 157651 257807 157699 257835
rect 157389 257773 157699 257807
rect 157389 257745 157437 257773
rect 157465 257745 157499 257773
rect 157527 257745 157561 257773
rect 157589 257745 157623 257773
rect 157651 257745 157699 257773
rect 157389 254075 157699 257745
rect 164529 299190 164839 299718
rect 164529 299162 164577 299190
rect 164605 299162 164639 299190
rect 164667 299162 164701 299190
rect 164729 299162 164763 299190
rect 164791 299162 164839 299190
rect 164529 299128 164839 299162
rect 164529 299100 164577 299128
rect 164605 299100 164639 299128
rect 164667 299100 164701 299128
rect 164729 299100 164763 299128
rect 164791 299100 164839 299128
rect 164529 299066 164839 299100
rect 164529 299038 164577 299066
rect 164605 299038 164639 299066
rect 164667 299038 164701 299066
rect 164729 299038 164763 299066
rect 164791 299038 164839 299066
rect 164529 299004 164839 299038
rect 164529 298976 164577 299004
rect 164605 298976 164639 299004
rect 164667 298976 164701 299004
rect 164729 298976 164763 299004
rect 164791 298976 164839 299004
rect 164529 290959 164839 298976
rect 164529 290931 164577 290959
rect 164605 290931 164639 290959
rect 164667 290931 164701 290959
rect 164729 290931 164763 290959
rect 164791 290931 164839 290959
rect 164529 290897 164839 290931
rect 164529 290869 164577 290897
rect 164605 290869 164639 290897
rect 164667 290869 164701 290897
rect 164729 290869 164763 290897
rect 164791 290869 164839 290897
rect 164529 290835 164839 290869
rect 164529 290807 164577 290835
rect 164605 290807 164639 290835
rect 164667 290807 164701 290835
rect 164729 290807 164763 290835
rect 164791 290807 164839 290835
rect 164529 290773 164839 290807
rect 164529 290745 164577 290773
rect 164605 290745 164639 290773
rect 164667 290745 164701 290773
rect 164729 290745 164763 290773
rect 164791 290745 164839 290773
rect 164529 281959 164839 290745
rect 164529 281931 164577 281959
rect 164605 281931 164639 281959
rect 164667 281931 164701 281959
rect 164729 281931 164763 281959
rect 164791 281931 164839 281959
rect 164529 281897 164839 281931
rect 164529 281869 164577 281897
rect 164605 281869 164639 281897
rect 164667 281869 164701 281897
rect 164729 281869 164763 281897
rect 164791 281869 164839 281897
rect 164529 281835 164839 281869
rect 164529 281807 164577 281835
rect 164605 281807 164639 281835
rect 164667 281807 164701 281835
rect 164729 281807 164763 281835
rect 164791 281807 164839 281835
rect 164529 281773 164839 281807
rect 164529 281745 164577 281773
rect 164605 281745 164639 281773
rect 164667 281745 164701 281773
rect 164729 281745 164763 281773
rect 164791 281745 164839 281773
rect 164529 272959 164839 281745
rect 164529 272931 164577 272959
rect 164605 272931 164639 272959
rect 164667 272931 164701 272959
rect 164729 272931 164763 272959
rect 164791 272931 164839 272959
rect 164529 272897 164839 272931
rect 164529 272869 164577 272897
rect 164605 272869 164639 272897
rect 164667 272869 164701 272897
rect 164729 272869 164763 272897
rect 164791 272869 164839 272897
rect 164529 272835 164839 272869
rect 164529 272807 164577 272835
rect 164605 272807 164639 272835
rect 164667 272807 164701 272835
rect 164729 272807 164763 272835
rect 164791 272807 164839 272835
rect 164529 272773 164839 272807
rect 164529 272745 164577 272773
rect 164605 272745 164639 272773
rect 164667 272745 164701 272773
rect 164729 272745 164763 272773
rect 164791 272745 164839 272773
rect 164529 263959 164839 272745
rect 164529 263931 164577 263959
rect 164605 263931 164639 263959
rect 164667 263931 164701 263959
rect 164729 263931 164763 263959
rect 164791 263931 164839 263959
rect 164529 263897 164839 263931
rect 164529 263869 164577 263897
rect 164605 263869 164639 263897
rect 164667 263869 164701 263897
rect 164729 263869 164763 263897
rect 164791 263869 164839 263897
rect 164529 263835 164839 263869
rect 164529 263807 164577 263835
rect 164605 263807 164639 263835
rect 164667 263807 164701 263835
rect 164729 263807 164763 263835
rect 164791 263807 164839 263835
rect 164529 263773 164839 263807
rect 164529 263745 164577 263773
rect 164605 263745 164639 263773
rect 164667 263745 164701 263773
rect 164729 263745 164763 263773
rect 164791 263745 164839 263773
rect 164529 254959 164839 263745
rect 164529 254931 164577 254959
rect 164605 254931 164639 254959
rect 164667 254931 164701 254959
rect 164729 254931 164763 254959
rect 164791 254931 164839 254959
rect 164529 254897 164839 254931
rect 164529 254869 164577 254897
rect 164605 254869 164639 254897
rect 164667 254869 164701 254897
rect 164729 254869 164763 254897
rect 164791 254869 164839 254897
rect 164529 254835 164839 254869
rect 164529 254807 164577 254835
rect 164605 254807 164639 254835
rect 164667 254807 164701 254835
rect 164729 254807 164763 254835
rect 164791 254807 164839 254835
rect 164529 254773 164839 254807
rect 164529 254745 164577 254773
rect 164605 254745 164639 254773
rect 164667 254745 164701 254773
rect 164729 254745 164763 254773
rect 164791 254745 164839 254773
rect 164529 254075 164839 254745
rect 166389 299670 166699 299718
rect 166389 299642 166437 299670
rect 166465 299642 166499 299670
rect 166527 299642 166561 299670
rect 166589 299642 166623 299670
rect 166651 299642 166699 299670
rect 166389 299608 166699 299642
rect 166389 299580 166437 299608
rect 166465 299580 166499 299608
rect 166527 299580 166561 299608
rect 166589 299580 166623 299608
rect 166651 299580 166699 299608
rect 166389 299546 166699 299580
rect 166389 299518 166437 299546
rect 166465 299518 166499 299546
rect 166527 299518 166561 299546
rect 166589 299518 166623 299546
rect 166651 299518 166699 299546
rect 166389 299484 166699 299518
rect 166389 299456 166437 299484
rect 166465 299456 166499 299484
rect 166527 299456 166561 299484
rect 166589 299456 166623 299484
rect 166651 299456 166699 299484
rect 166389 293959 166699 299456
rect 166389 293931 166437 293959
rect 166465 293931 166499 293959
rect 166527 293931 166561 293959
rect 166589 293931 166623 293959
rect 166651 293931 166699 293959
rect 166389 293897 166699 293931
rect 166389 293869 166437 293897
rect 166465 293869 166499 293897
rect 166527 293869 166561 293897
rect 166589 293869 166623 293897
rect 166651 293869 166699 293897
rect 166389 293835 166699 293869
rect 166389 293807 166437 293835
rect 166465 293807 166499 293835
rect 166527 293807 166561 293835
rect 166589 293807 166623 293835
rect 166651 293807 166699 293835
rect 166389 293773 166699 293807
rect 166389 293745 166437 293773
rect 166465 293745 166499 293773
rect 166527 293745 166561 293773
rect 166589 293745 166623 293773
rect 166651 293745 166699 293773
rect 166389 284959 166699 293745
rect 166389 284931 166437 284959
rect 166465 284931 166499 284959
rect 166527 284931 166561 284959
rect 166589 284931 166623 284959
rect 166651 284931 166699 284959
rect 166389 284897 166699 284931
rect 166389 284869 166437 284897
rect 166465 284869 166499 284897
rect 166527 284869 166561 284897
rect 166589 284869 166623 284897
rect 166651 284869 166699 284897
rect 166389 284835 166699 284869
rect 166389 284807 166437 284835
rect 166465 284807 166499 284835
rect 166527 284807 166561 284835
rect 166589 284807 166623 284835
rect 166651 284807 166699 284835
rect 166389 284773 166699 284807
rect 166389 284745 166437 284773
rect 166465 284745 166499 284773
rect 166527 284745 166561 284773
rect 166589 284745 166623 284773
rect 166651 284745 166699 284773
rect 166389 275959 166699 284745
rect 166389 275931 166437 275959
rect 166465 275931 166499 275959
rect 166527 275931 166561 275959
rect 166589 275931 166623 275959
rect 166651 275931 166699 275959
rect 166389 275897 166699 275931
rect 166389 275869 166437 275897
rect 166465 275869 166499 275897
rect 166527 275869 166561 275897
rect 166589 275869 166623 275897
rect 166651 275869 166699 275897
rect 166389 275835 166699 275869
rect 166389 275807 166437 275835
rect 166465 275807 166499 275835
rect 166527 275807 166561 275835
rect 166589 275807 166623 275835
rect 166651 275807 166699 275835
rect 166389 275773 166699 275807
rect 166389 275745 166437 275773
rect 166465 275745 166499 275773
rect 166527 275745 166561 275773
rect 166589 275745 166623 275773
rect 166651 275745 166699 275773
rect 166389 266959 166699 275745
rect 166389 266931 166437 266959
rect 166465 266931 166499 266959
rect 166527 266931 166561 266959
rect 166589 266931 166623 266959
rect 166651 266931 166699 266959
rect 166389 266897 166699 266931
rect 166389 266869 166437 266897
rect 166465 266869 166499 266897
rect 166527 266869 166561 266897
rect 166589 266869 166623 266897
rect 166651 266869 166699 266897
rect 166389 266835 166699 266869
rect 166389 266807 166437 266835
rect 166465 266807 166499 266835
rect 166527 266807 166561 266835
rect 166589 266807 166623 266835
rect 166651 266807 166699 266835
rect 166389 266773 166699 266807
rect 166389 266745 166437 266773
rect 166465 266745 166499 266773
rect 166527 266745 166561 266773
rect 166589 266745 166623 266773
rect 166651 266745 166699 266773
rect 166389 257959 166699 266745
rect 166389 257931 166437 257959
rect 166465 257931 166499 257959
rect 166527 257931 166561 257959
rect 166589 257931 166623 257959
rect 166651 257931 166699 257959
rect 166389 257897 166699 257931
rect 166389 257869 166437 257897
rect 166465 257869 166499 257897
rect 166527 257869 166561 257897
rect 166589 257869 166623 257897
rect 166651 257869 166699 257897
rect 166389 257835 166699 257869
rect 166389 257807 166437 257835
rect 166465 257807 166499 257835
rect 166527 257807 166561 257835
rect 166589 257807 166623 257835
rect 166651 257807 166699 257835
rect 166389 257773 166699 257807
rect 166389 257745 166437 257773
rect 166465 257745 166499 257773
rect 166527 257745 166561 257773
rect 166589 257745 166623 257773
rect 166651 257745 166699 257773
rect 166389 254075 166699 257745
rect 173529 299190 173839 299718
rect 173529 299162 173577 299190
rect 173605 299162 173639 299190
rect 173667 299162 173701 299190
rect 173729 299162 173763 299190
rect 173791 299162 173839 299190
rect 173529 299128 173839 299162
rect 173529 299100 173577 299128
rect 173605 299100 173639 299128
rect 173667 299100 173701 299128
rect 173729 299100 173763 299128
rect 173791 299100 173839 299128
rect 173529 299066 173839 299100
rect 173529 299038 173577 299066
rect 173605 299038 173639 299066
rect 173667 299038 173701 299066
rect 173729 299038 173763 299066
rect 173791 299038 173839 299066
rect 173529 299004 173839 299038
rect 173529 298976 173577 299004
rect 173605 298976 173639 299004
rect 173667 298976 173701 299004
rect 173729 298976 173763 299004
rect 173791 298976 173839 299004
rect 173529 290959 173839 298976
rect 173529 290931 173577 290959
rect 173605 290931 173639 290959
rect 173667 290931 173701 290959
rect 173729 290931 173763 290959
rect 173791 290931 173839 290959
rect 173529 290897 173839 290931
rect 173529 290869 173577 290897
rect 173605 290869 173639 290897
rect 173667 290869 173701 290897
rect 173729 290869 173763 290897
rect 173791 290869 173839 290897
rect 173529 290835 173839 290869
rect 173529 290807 173577 290835
rect 173605 290807 173639 290835
rect 173667 290807 173701 290835
rect 173729 290807 173763 290835
rect 173791 290807 173839 290835
rect 173529 290773 173839 290807
rect 173529 290745 173577 290773
rect 173605 290745 173639 290773
rect 173667 290745 173701 290773
rect 173729 290745 173763 290773
rect 173791 290745 173839 290773
rect 173529 281959 173839 290745
rect 173529 281931 173577 281959
rect 173605 281931 173639 281959
rect 173667 281931 173701 281959
rect 173729 281931 173763 281959
rect 173791 281931 173839 281959
rect 173529 281897 173839 281931
rect 173529 281869 173577 281897
rect 173605 281869 173639 281897
rect 173667 281869 173701 281897
rect 173729 281869 173763 281897
rect 173791 281869 173839 281897
rect 173529 281835 173839 281869
rect 173529 281807 173577 281835
rect 173605 281807 173639 281835
rect 173667 281807 173701 281835
rect 173729 281807 173763 281835
rect 173791 281807 173839 281835
rect 173529 281773 173839 281807
rect 173529 281745 173577 281773
rect 173605 281745 173639 281773
rect 173667 281745 173701 281773
rect 173729 281745 173763 281773
rect 173791 281745 173839 281773
rect 173529 272959 173839 281745
rect 173529 272931 173577 272959
rect 173605 272931 173639 272959
rect 173667 272931 173701 272959
rect 173729 272931 173763 272959
rect 173791 272931 173839 272959
rect 173529 272897 173839 272931
rect 173529 272869 173577 272897
rect 173605 272869 173639 272897
rect 173667 272869 173701 272897
rect 173729 272869 173763 272897
rect 173791 272869 173839 272897
rect 173529 272835 173839 272869
rect 173529 272807 173577 272835
rect 173605 272807 173639 272835
rect 173667 272807 173701 272835
rect 173729 272807 173763 272835
rect 173791 272807 173839 272835
rect 173529 272773 173839 272807
rect 173529 272745 173577 272773
rect 173605 272745 173639 272773
rect 173667 272745 173701 272773
rect 173729 272745 173763 272773
rect 173791 272745 173839 272773
rect 173529 263959 173839 272745
rect 173529 263931 173577 263959
rect 173605 263931 173639 263959
rect 173667 263931 173701 263959
rect 173729 263931 173763 263959
rect 173791 263931 173839 263959
rect 173529 263897 173839 263931
rect 173529 263869 173577 263897
rect 173605 263869 173639 263897
rect 173667 263869 173701 263897
rect 173729 263869 173763 263897
rect 173791 263869 173839 263897
rect 173529 263835 173839 263869
rect 173529 263807 173577 263835
rect 173605 263807 173639 263835
rect 173667 263807 173701 263835
rect 173729 263807 173763 263835
rect 173791 263807 173839 263835
rect 173529 263773 173839 263807
rect 173529 263745 173577 263773
rect 173605 263745 173639 263773
rect 173667 263745 173701 263773
rect 173729 263745 173763 263773
rect 173791 263745 173839 263773
rect 173529 254959 173839 263745
rect 173529 254931 173577 254959
rect 173605 254931 173639 254959
rect 173667 254931 173701 254959
rect 173729 254931 173763 254959
rect 173791 254931 173839 254959
rect 173529 254897 173839 254931
rect 173529 254869 173577 254897
rect 173605 254869 173639 254897
rect 173667 254869 173701 254897
rect 173729 254869 173763 254897
rect 173791 254869 173839 254897
rect 173529 254835 173839 254869
rect 173529 254807 173577 254835
rect 173605 254807 173639 254835
rect 173667 254807 173701 254835
rect 173729 254807 173763 254835
rect 173791 254807 173839 254835
rect 173529 254773 173839 254807
rect 173529 254745 173577 254773
rect 173605 254745 173639 254773
rect 173667 254745 173701 254773
rect 173729 254745 173763 254773
rect 173791 254745 173839 254773
rect 173529 254075 173839 254745
rect 175389 299670 175699 299718
rect 175389 299642 175437 299670
rect 175465 299642 175499 299670
rect 175527 299642 175561 299670
rect 175589 299642 175623 299670
rect 175651 299642 175699 299670
rect 175389 299608 175699 299642
rect 175389 299580 175437 299608
rect 175465 299580 175499 299608
rect 175527 299580 175561 299608
rect 175589 299580 175623 299608
rect 175651 299580 175699 299608
rect 175389 299546 175699 299580
rect 175389 299518 175437 299546
rect 175465 299518 175499 299546
rect 175527 299518 175561 299546
rect 175589 299518 175623 299546
rect 175651 299518 175699 299546
rect 175389 299484 175699 299518
rect 175389 299456 175437 299484
rect 175465 299456 175499 299484
rect 175527 299456 175561 299484
rect 175589 299456 175623 299484
rect 175651 299456 175699 299484
rect 175389 293959 175699 299456
rect 175389 293931 175437 293959
rect 175465 293931 175499 293959
rect 175527 293931 175561 293959
rect 175589 293931 175623 293959
rect 175651 293931 175699 293959
rect 175389 293897 175699 293931
rect 175389 293869 175437 293897
rect 175465 293869 175499 293897
rect 175527 293869 175561 293897
rect 175589 293869 175623 293897
rect 175651 293869 175699 293897
rect 175389 293835 175699 293869
rect 175389 293807 175437 293835
rect 175465 293807 175499 293835
rect 175527 293807 175561 293835
rect 175589 293807 175623 293835
rect 175651 293807 175699 293835
rect 175389 293773 175699 293807
rect 175389 293745 175437 293773
rect 175465 293745 175499 293773
rect 175527 293745 175561 293773
rect 175589 293745 175623 293773
rect 175651 293745 175699 293773
rect 175389 284959 175699 293745
rect 175389 284931 175437 284959
rect 175465 284931 175499 284959
rect 175527 284931 175561 284959
rect 175589 284931 175623 284959
rect 175651 284931 175699 284959
rect 175389 284897 175699 284931
rect 175389 284869 175437 284897
rect 175465 284869 175499 284897
rect 175527 284869 175561 284897
rect 175589 284869 175623 284897
rect 175651 284869 175699 284897
rect 175389 284835 175699 284869
rect 175389 284807 175437 284835
rect 175465 284807 175499 284835
rect 175527 284807 175561 284835
rect 175589 284807 175623 284835
rect 175651 284807 175699 284835
rect 175389 284773 175699 284807
rect 175389 284745 175437 284773
rect 175465 284745 175499 284773
rect 175527 284745 175561 284773
rect 175589 284745 175623 284773
rect 175651 284745 175699 284773
rect 175389 275959 175699 284745
rect 175389 275931 175437 275959
rect 175465 275931 175499 275959
rect 175527 275931 175561 275959
rect 175589 275931 175623 275959
rect 175651 275931 175699 275959
rect 175389 275897 175699 275931
rect 175389 275869 175437 275897
rect 175465 275869 175499 275897
rect 175527 275869 175561 275897
rect 175589 275869 175623 275897
rect 175651 275869 175699 275897
rect 175389 275835 175699 275869
rect 175389 275807 175437 275835
rect 175465 275807 175499 275835
rect 175527 275807 175561 275835
rect 175589 275807 175623 275835
rect 175651 275807 175699 275835
rect 175389 275773 175699 275807
rect 175389 275745 175437 275773
rect 175465 275745 175499 275773
rect 175527 275745 175561 275773
rect 175589 275745 175623 275773
rect 175651 275745 175699 275773
rect 175389 266959 175699 275745
rect 175389 266931 175437 266959
rect 175465 266931 175499 266959
rect 175527 266931 175561 266959
rect 175589 266931 175623 266959
rect 175651 266931 175699 266959
rect 175389 266897 175699 266931
rect 175389 266869 175437 266897
rect 175465 266869 175499 266897
rect 175527 266869 175561 266897
rect 175589 266869 175623 266897
rect 175651 266869 175699 266897
rect 175389 266835 175699 266869
rect 175389 266807 175437 266835
rect 175465 266807 175499 266835
rect 175527 266807 175561 266835
rect 175589 266807 175623 266835
rect 175651 266807 175699 266835
rect 175389 266773 175699 266807
rect 175389 266745 175437 266773
rect 175465 266745 175499 266773
rect 175527 266745 175561 266773
rect 175589 266745 175623 266773
rect 175651 266745 175699 266773
rect 175389 257959 175699 266745
rect 175389 257931 175437 257959
rect 175465 257931 175499 257959
rect 175527 257931 175561 257959
rect 175589 257931 175623 257959
rect 175651 257931 175699 257959
rect 175389 257897 175699 257931
rect 175389 257869 175437 257897
rect 175465 257869 175499 257897
rect 175527 257869 175561 257897
rect 175589 257869 175623 257897
rect 175651 257869 175699 257897
rect 175389 257835 175699 257869
rect 175389 257807 175437 257835
rect 175465 257807 175499 257835
rect 175527 257807 175561 257835
rect 175589 257807 175623 257835
rect 175651 257807 175699 257835
rect 175389 257773 175699 257807
rect 175389 257745 175437 257773
rect 175465 257745 175499 257773
rect 175527 257745 175561 257773
rect 175589 257745 175623 257773
rect 175651 257745 175699 257773
rect 175389 254075 175699 257745
rect 182529 299190 182839 299718
rect 182529 299162 182577 299190
rect 182605 299162 182639 299190
rect 182667 299162 182701 299190
rect 182729 299162 182763 299190
rect 182791 299162 182839 299190
rect 182529 299128 182839 299162
rect 182529 299100 182577 299128
rect 182605 299100 182639 299128
rect 182667 299100 182701 299128
rect 182729 299100 182763 299128
rect 182791 299100 182839 299128
rect 182529 299066 182839 299100
rect 182529 299038 182577 299066
rect 182605 299038 182639 299066
rect 182667 299038 182701 299066
rect 182729 299038 182763 299066
rect 182791 299038 182839 299066
rect 182529 299004 182839 299038
rect 182529 298976 182577 299004
rect 182605 298976 182639 299004
rect 182667 298976 182701 299004
rect 182729 298976 182763 299004
rect 182791 298976 182839 299004
rect 182529 290959 182839 298976
rect 182529 290931 182577 290959
rect 182605 290931 182639 290959
rect 182667 290931 182701 290959
rect 182729 290931 182763 290959
rect 182791 290931 182839 290959
rect 182529 290897 182839 290931
rect 182529 290869 182577 290897
rect 182605 290869 182639 290897
rect 182667 290869 182701 290897
rect 182729 290869 182763 290897
rect 182791 290869 182839 290897
rect 182529 290835 182839 290869
rect 182529 290807 182577 290835
rect 182605 290807 182639 290835
rect 182667 290807 182701 290835
rect 182729 290807 182763 290835
rect 182791 290807 182839 290835
rect 182529 290773 182839 290807
rect 182529 290745 182577 290773
rect 182605 290745 182639 290773
rect 182667 290745 182701 290773
rect 182729 290745 182763 290773
rect 182791 290745 182839 290773
rect 182529 281959 182839 290745
rect 182529 281931 182577 281959
rect 182605 281931 182639 281959
rect 182667 281931 182701 281959
rect 182729 281931 182763 281959
rect 182791 281931 182839 281959
rect 182529 281897 182839 281931
rect 182529 281869 182577 281897
rect 182605 281869 182639 281897
rect 182667 281869 182701 281897
rect 182729 281869 182763 281897
rect 182791 281869 182839 281897
rect 182529 281835 182839 281869
rect 182529 281807 182577 281835
rect 182605 281807 182639 281835
rect 182667 281807 182701 281835
rect 182729 281807 182763 281835
rect 182791 281807 182839 281835
rect 182529 281773 182839 281807
rect 182529 281745 182577 281773
rect 182605 281745 182639 281773
rect 182667 281745 182701 281773
rect 182729 281745 182763 281773
rect 182791 281745 182839 281773
rect 182529 272959 182839 281745
rect 182529 272931 182577 272959
rect 182605 272931 182639 272959
rect 182667 272931 182701 272959
rect 182729 272931 182763 272959
rect 182791 272931 182839 272959
rect 182529 272897 182839 272931
rect 182529 272869 182577 272897
rect 182605 272869 182639 272897
rect 182667 272869 182701 272897
rect 182729 272869 182763 272897
rect 182791 272869 182839 272897
rect 182529 272835 182839 272869
rect 182529 272807 182577 272835
rect 182605 272807 182639 272835
rect 182667 272807 182701 272835
rect 182729 272807 182763 272835
rect 182791 272807 182839 272835
rect 182529 272773 182839 272807
rect 182529 272745 182577 272773
rect 182605 272745 182639 272773
rect 182667 272745 182701 272773
rect 182729 272745 182763 272773
rect 182791 272745 182839 272773
rect 182529 263959 182839 272745
rect 182529 263931 182577 263959
rect 182605 263931 182639 263959
rect 182667 263931 182701 263959
rect 182729 263931 182763 263959
rect 182791 263931 182839 263959
rect 182529 263897 182839 263931
rect 182529 263869 182577 263897
rect 182605 263869 182639 263897
rect 182667 263869 182701 263897
rect 182729 263869 182763 263897
rect 182791 263869 182839 263897
rect 182529 263835 182839 263869
rect 182529 263807 182577 263835
rect 182605 263807 182639 263835
rect 182667 263807 182701 263835
rect 182729 263807 182763 263835
rect 182791 263807 182839 263835
rect 182529 263773 182839 263807
rect 182529 263745 182577 263773
rect 182605 263745 182639 263773
rect 182667 263745 182701 263773
rect 182729 263745 182763 263773
rect 182791 263745 182839 263773
rect 182529 254959 182839 263745
rect 182529 254931 182577 254959
rect 182605 254931 182639 254959
rect 182667 254931 182701 254959
rect 182729 254931 182763 254959
rect 182791 254931 182839 254959
rect 182529 254897 182839 254931
rect 182529 254869 182577 254897
rect 182605 254869 182639 254897
rect 182667 254869 182701 254897
rect 182729 254869 182763 254897
rect 182791 254869 182839 254897
rect 182529 254835 182839 254869
rect 182529 254807 182577 254835
rect 182605 254807 182639 254835
rect 182667 254807 182701 254835
rect 182729 254807 182763 254835
rect 182791 254807 182839 254835
rect 182529 254773 182839 254807
rect 182529 254745 182577 254773
rect 182605 254745 182639 254773
rect 182667 254745 182701 254773
rect 182729 254745 182763 254773
rect 182791 254745 182839 254773
rect 182529 254075 182839 254745
rect 184389 299670 184699 299718
rect 184389 299642 184437 299670
rect 184465 299642 184499 299670
rect 184527 299642 184561 299670
rect 184589 299642 184623 299670
rect 184651 299642 184699 299670
rect 184389 299608 184699 299642
rect 184389 299580 184437 299608
rect 184465 299580 184499 299608
rect 184527 299580 184561 299608
rect 184589 299580 184623 299608
rect 184651 299580 184699 299608
rect 184389 299546 184699 299580
rect 184389 299518 184437 299546
rect 184465 299518 184499 299546
rect 184527 299518 184561 299546
rect 184589 299518 184623 299546
rect 184651 299518 184699 299546
rect 184389 299484 184699 299518
rect 184389 299456 184437 299484
rect 184465 299456 184499 299484
rect 184527 299456 184561 299484
rect 184589 299456 184623 299484
rect 184651 299456 184699 299484
rect 184389 293959 184699 299456
rect 184389 293931 184437 293959
rect 184465 293931 184499 293959
rect 184527 293931 184561 293959
rect 184589 293931 184623 293959
rect 184651 293931 184699 293959
rect 184389 293897 184699 293931
rect 184389 293869 184437 293897
rect 184465 293869 184499 293897
rect 184527 293869 184561 293897
rect 184589 293869 184623 293897
rect 184651 293869 184699 293897
rect 184389 293835 184699 293869
rect 184389 293807 184437 293835
rect 184465 293807 184499 293835
rect 184527 293807 184561 293835
rect 184589 293807 184623 293835
rect 184651 293807 184699 293835
rect 184389 293773 184699 293807
rect 184389 293745 184437 293773
rect 184465 293745 184499 293773
rect 184527 293745 184561 293773
rect 184589 293745 184623 293773
rect 184651 293745 184699 293773
rect 184389 284959 184699 293745
rect 184389 284931 184437 284959
rect 184465 284931 184499 284959
rect 184527 284931 184561 284959
rect 184589 284931 184623 284959
rect 184651 284931 184699 284959
rect 184389 284897 184699 284931
rect 184389 284869 184437 284897
rect 184465 284869 184499 284897
rect 184527 284869 184561 284897
rect 184589 284869 184623 284897
rect 184651 284869 184699 284897
rect 184389 284835 184699 284869
rect 184389 284807 184437 284835
rect 184465 284807 184499 284835
rect 184527 284807 184561 284835
rect 184589 284807 184623 284835
rect 184651 284807 184699 284835
rect 184389 284773 184699 284807
rect 184389 284745 184437 284773
rect 184465 284745 184499 284773
rect 184527 284745 184561 284773
rect 184589 284745 184623 284773
rect 184651 284745 184699 284773
rect 184389 275959 184699 284745
rect 184389 275931 184437 275959
rect 184465 275931 184499 275959
rect 184527 275931 184561 275959
rect 184589 275931 184623 275959
rect 184651 275931 184699 275959
rect 184389 275897 184699 275931
rect 184389 275869 184437 275897
rect 184465 275869 184499 275897
rect 184527 275869 184561 275897
rect 184589 275869 184623 275897
rect 184651 275869 184699 275897
rect 184389 275835 184699 275869
rect 184389 275807 184437 275835
rect 184465 275807 184499 275835
rect 184527 275807 184561 275835
rect 184589 275807 184623 275835
rect 184651 275807 184699 275835
rect 184389 275773 184699 275807
rect 184389 275745 184437 275773
rect 184465 275745 184499 275773
rect 184527 275745 184561 275773
rect 184589 275745 184623 275773
rect 184651 275745 184699 275773
rect 184389 266959 184699 275745
rect 184389 266931 184437 266959
rect 184465 266931 184499 266959
rect 184527 266931 184561 266959
rect 184589 266931 184623 266959
rect 184651 266931 184699 266959
rect 184389 266897 184699 266931
rect 184389 266869 184437 266897
rect 184465 266869 184499 266897
rect 184527 266869 184561 266897
rect 184589 266869 184623 266897
rect 184651 266869 184699 266897
rect 184389 266835 184699 266869
rect 184389 266807 184437 266835
rect 184465 266807 184499 266835
rect 184527 266807 184561 266835
rect 184589 266807 184623 266835
rect 184651 266807 184699 266835
rect 184389 266773 184699 266807
rect 184389 266745 184437 266773
rect 184465 266745 184499 266773
rect 184527 266745 184561 266773
rect 184589 266745 184623 266773
rect 184651 266745 184699 266773
rect 184389 257959 184699 266745
rect 184389 257931 184437 257959
rect 184465 257931 184499 257959
rect 184527 257931 184561 257959
rect 184589 257931 184623 257959
rect 184651 257931 184699 257959
rect 184389 257897 184699 257931
rect 184389 257869 184437 257897
rect 184465 257869 184499 257897
rect 184527 257869 184561 257897
rect 184589 257869 184623 257897
rect 184651 257869 184699 257897
rect 184389 257835 184699 257869
rect 184389 257807 184437 257835
rect 184465 257807 184499 257835
rect 184527 257807 184561 257835
rect 184589 257807 184623 257835
rect 184651 257807 184699 257835
rect 184389 257773 184699 257807
rect 184389 257745 184437 257773
rect 184465 257745 184499 257773
rect 184527 257745 184561 257773
rect 184589 257745 184623 257773
rect 184651 257745 184699 257773
rect 184389 254075 184699 257745
rect 191529 299190 191839 299718
rect 191529 299162 191577 299190
rect 191605 299162 191639 299190
rect 191667 299162 191701 299190
rect 191729 299162 191763 299190
rect 191791 299162 191839 299190
rect 191529 299128 191839 299162
rect 191529 299100 191577 299128
rect 191605 299100 191639 299128
rect 191667 299100 191701 299128
rect 191729 299100 191763 299128
rect 191791 299100 191839 299128
rect 191529 299066 191839 299100
rect 191529 299038 191577 299066
rect 191605 299038 191639 299066
rect 191667 299038 191701 299066
rect 191729 299038 191763 299066
rect 191791 299038 191839 299066
rect 191529 299004 191839 299038
rect 191529 298976 191577 299004
rect 191605 298976 191639 299004
rect 191667 298976 191701 299004
rect 191729 298976 191763 299004
rect 191791 298976 191839 299004
rect 191529 290959 191839 298976
rect 191529 290931 191577 290959
rect 191605 290931 191639 290959
rect 191667 290931 191701 290959
rect 191729 290931 191763 290959
rect 191791 290931 191839 290959
rect 191529 290897 191839 290931
rect 191529 290869 191577 290897
rect 191605 290869 191639 290897
rect 191667 290869 191701 290897
rect 191729 290869 191763 290897
rect 191791 290869 191839 290897
rect 191529 290835 191839 290869
rect 191529 290807 191577 290835
rect 191605 290807 191639 290835
rect 191667 290807 191701 290835
rect 191729 290807 191763 290835
rect 191791 290807 191839 290835
rect 191529 290773 191839 290807
rect 191529 290745 191577 290773
rect 191605 290745 191639 290773
rect 191667 290745 191701 290773
rect 191729 290745 191763 290773
rect 191791 290745 191839 290773
rect 191529 281959 191839 290745
rect 191529 281931 191577 281959
rect 191605 281931 191639 281959
rect 191667 281931 191701 281959
rect 191729 281931 191763 281959
rect 191791 281931 191839 281959
rect 191529 281897 191839 281931
rect 191529 281869 191577 281897
rect 191605 281869 191639 281897
rect 191667 281869 191701 281897
rect 191729 281869 191763 281897
rect 191791 281869 191839 281897
rect 191529 281835 191839 281869
rect 191529 281807 191577 281835
rect 191605 281807 191639 281835
rect 191667 281807 191701 281835
rect 191729 281807 191763 281835
rect 191791 281807 191839 281835
rect 191529 281773 191839 281807
rect 191529 281745 191577 281773
rect 191605 281745 191639 281773
rect 191667 281745 191701 281773
rect 191729 281745 191763 281773
rect 191791 281745 191839 281773
rect 191529 272959 191839 281745
rect 191529 272931 191577 272959
rect 191605 272931 191639 272959
rect 191667 272931 191701 272959
rect 191729 272931 191763 272959
rect 191791 272931 191839 272959
rect 191529 272897 191839 272931
rect 191529 272869 191577 272897
rect 191605 272869 191639 272897
rect 191667 272869 191701 272897
rect 191729 272869 191763 272897
rect 191791 272869 191839 272897
rect 191529 272835 191839 272869
rect 191529 272807 191577 272835
rect 191605 272807 191639 272835
rect 191667 272807 191701 272835
rect 191729 272807 191763 272835
rect 191791 272807 191839 272835
rect 191529 272773 191839 272807
rect 191529 272745 191577 272773
rect 191605 272745 191639 272773
rect 191667 272745 191701 272773
rect 191729 272745 191763 272773
rect 191791 272745 191839 272773
rect 191529 263959 191839 272745
rect 191529 263931 191577 263959
rect 191605 263931 191639 263959
rect 191667 263931 191701 263959
rect 191729 263931 191763 263959
rect 191791 263931 191839 263959
rect 191529 263897 191839 263931
rect 191529 263869 191577 263897
rect 191605 263869 191639 263897
rect 191667 263869 191701 263897
rect 191729 263869 191763 263897
rect 191791 263869 191839 263897
rect 191529 263835 191839 263869
rect 191529 263807 191577 263835
rect 191605 263807 191639 263835
rect 191667 263807 191701 263835
rect 191729 263807 191763 263835
rect 191791 263807 191839 263835
rect 191529 263773 191839 263807
rect 191529 263745 191577 263773
rect 191605 263745 191639 263773
rect 191667 263745 191701 263773
rect 191729 263745 191763 263773
rect 191791 263745 191839 263773
rect 191529 254959 191839 263745
rect 191529 254931 191577 254959
rect 191605 254931 191639 254959
rect 191667 254931 191701 254959
rect 191729 254931 191763 254959
rect 191791 254931 191839 254959
rect 191529 254897 191839 254931
rect 191529 254869 191577 254897
rect 191605 254869 191639 254897
rect 191667 254869 191701 254897
rect 191729 254869 191763 254897
rect 191791 254869 191839 254897
rect 191529 254835 191839 254869
rect 191529 254807 191577 254835
rect 191605 254807 191639 254835
rect 191667 254807 191701 254835
rect 191729 254807 191763 254835
rect 191791 254807 191839 254835
rect 191529 254773 191839 254807
rect 191529 254745 191577 254773
rect 191605 254745 191639 254773
rect 191667 254745 191701 254773
rect 191729 254745 191763 254773
rect 191791 254745 191839 254773
rect 191529 254075 191839 254745
rect 193389 299670 193699 299718
rect 193389 299642 193437 299670
rect 193465 299642 193499 299670
rect 193527 299642 193561 299670
rect 193589 299642 193623 299670
rect 193651 299642 193699 299670
rect 193389 299608 193699 299642
rect 193389 299580 193437 299608
rect 193465 299580 193499 299608
rect 193527 299580 193561 299608
rect 193589 299580 193623 299608
rect 193651 299580 193699 299608
rect 193389 299546 193699 299580
rect 193389 299518 193437 299546
rect 193465 299518 193499 299546
rect 193527 299518 193561 299546
rect 193589 299518 193623 299546
rect 193651 299518 193699 299546
rect 193389 299484 193699 299518
rect 193389 299456 193437 299484
rect 193465 299456 193499 299484
rect 193527 299456 193561 299484
rect 193589 299456 193623 299484
rect 193651 299456 193699 299484
rect 193389 293959 193699 299456
rect 193389 293931 193437 293959
rect 193465 293931 193499 293959
rect 193527 293931 193561 293959
rect 193589 293931 193623 293959
rect 193651 293931 193699 293959
rect 193389 293897 193699 293931
rect 193389 293869 193437 293897
rect 193465 293869 193499 293897
rect 193527 293869 193561 293897
rect 193589 293869 193623 293897
rect 193651 293869 193699 293897
rect 193389 293835 193699 293869
rect 193389 293807 193437 293835
rect 193465 293807 193499 293835
rect 193527 293807 193561 293835
rect 193589 293807 193623 293835
rect 193651 293807 193699 293835
rect 193389 293773 193699 293807
rect 193389 293745 193437 293773
rect 193465 293745 193499 293773
rect 193527 293745 193561 293773
rect 193589 293745 193623 293773
rect 193651 293745 193699 293773
rect 193389 284959 193699 293745
rect 193389 284931 193437 284959
rect 193465 284931 193499 284959
rect 193527 284931 193561 284959
rect 193589 284931 193623 284959
rect 193651 284931 193699 284959
rect 193389 284897 193699 284931
rect 193389 284869 193437 284897
rect 193465 284869 193499 284897
rect 193527 284869 193561 284897
rect 193589 284869 193623 284897
rect 193651 284869 193699 284897
rect 193389 284835 193699 284869
rect 193389 284807 193437 284835
rect 193465 284807 193499 284835
rect 193527 284807 193561 284835
rect 193589 284807 193623 284835
rect 193651 284807 193699 284835
rect 193389 284773 193699 284807
rect 193389 284745 193437 284773
rect 193465 284745 193499 284773
rect 193527 284745 193561 284773
rect 193589 284745 193623 284773
rect 193651 284745 193699 284773
rect 193389 275959 193699 284745
rect 193389 275931 193437 275959
rect 193465 275931 193499 275959
rect 193527 275931 193561 275959
rect 193589 275931 193623 275959
rect 193651 275931 193699 275959
rect 193389 275897 193699 275931
rect 193389 275869 193437 275897
rect 193465 275869 193499 275897
rect 193527 275869 193561 275897
rect 193589 275869 193623 275897
rect 193651 275869 193699 275897
rect 193389 275835 193699 275869
rect 193389 275807 193437 275835
rect 193465 275807 193499 275835
rect 193527 275807 193561 275835
rect 193589 275807 193623 275835
rect 193651 275807 193699 275835
rect 193389 275773 193699 275807
rect 193389 275745 193437 275773
rect 193465 275745 193499 275773
rect 193527 275745 193561 275773
rect 193589 275745 193623 275773
rect 193651 275745 193699 275773
rect 193389 266959 193699 275745
rect 193389 266931 193437 266959
rect 193465 266931 193499 266959
rect 193527 266931 193561 266959
rect 193589 266931 193623 266959
rect 193651 266931 193699 266959
rect 193389 266897 193699 266931
rect 193389 266869 193437 266897
rect 193465 266869 193499 266897
rect 193527 266869 193561 266897
rect 193589 266869 193623 266897
rect 193651 266869 193699 266897
rect 193389 266835 193699 266869
rect 193389 266807 193437 266835
rect 193465 266807 193499 266835
rect 193527 266807 193561 266835
rect 193589 266807 193623 266835
rect 193651 266807 193699 266835
rect 193389 266773 193699 266807
rect 193389 266745 193437 266773
rect 193465 266745 193499 266773
rect 193527 266745 193561 266773
rect 193589 266745 193623 266773
rect 193651 266745 193699 266773
rect 193389 257959 193699 266745
rect 193389 257931 193437 257959
rect 193465 257931 193499 257959
rect 193527 257931 193561 257959
rect 193589 257931 193623 257959
rect 193651 257931 193699 257959
rect 193389 257897 193699 257931
rect 193389 257869 193437 257897
rect 193465 257869 193499 257897
rect 193527 257869 193561 257897
rect 193589 257869 193623 257897
rect 193651 257869 193699 257897
rect 193389 257835 193699 257869
rect 193389 257807 193437 257835
rect 193465 257807 193499 257835
rect 193527 257807 193561 257835
rect 193589 257807 193623 257835
rect 193651 257807 193699 257835
rect 193389 257773 193699 257807
rect 193389 257745 193437 257773
rect 193465 257745 193499 257773
rect 193527 257745 193561 257773
rect 193589 257745 193623 257773
rect 193651 257745 193699 257773
rect 193389 254075 193699 257745
rect 200529 299190 200839 299718
rect 200529 299162 200577 299190
rect 200605 299162 200639 299190
rect 200667 299162 200701 299190
rect 200729 299162 200763 299190
rect 200791 299162 200839 299190
rect 200529 299128 200839 299162
rect 200529 299100 200577 299128
rect 200605 299100 200639 299128
rect 200667 299100 200701 299128
rect 200729 299100 200763 299128
rect 200791 299100 200839 299128
rect 200529 299066 200839 299100
rect 200529 299038 200577 299066
rect 200605 299038 200639 299066
rect 200667 299038 200701 299066
rect 200729 299038 200763 299066
rect 200791 299038 200839 299066
rect 200529 299004 200839 299038
rect 200529 298976 200577 299004
rect 200605 298976 200639 299004
rect 200667 298976 200701 299004
rect 200729 298976 200763 299004
rect 200791 298976 200839 299004
rect 200529 290959 200839 298976
rect 200529 290931 200577 290959
rect 200605 290931 200639 290959
rect 200667 290931 200701 290959
rect 200729 290931 200763 290959
rect 200791 290931 200839 290959
rect 200529 290897 200839 290931
rect 200529 290869 200577 290897
rect 200605 290869 200639 290897
rect 200667 290869 200701 290897
rect 200729 290869 200763 290897
rect 200791 290869 200839 290897
rect 200529 290835 200839 290869
rect 200529 290807 200577 290835
rect 200605 290807 200639 290835
rect 200667 290807 200701 290835
rect 200729 290807 200763 290835
rect 200791 290807 200839 290835
rect 200529 290773 200839 290807
rect 200529 290745 200577 290773
rect 200605 290745 200639 290773
rect 200667 290745 200701 290773
rect 200729 290745 200763 290773
rect 200791 290745 200839 290773
rect 200529 281959 200839 290745
rect 200529 281931 200577 281959
rect 200605 281931 200639 281959
rect 200667 281931 200701 281959
rect 200729 281931 200763 281959
rect 200791 281931 200839 281959
rect 200529 281897 200839 281931
rect 200529 281869 200577 281897
rect 200605 281869 200639 281897
rect 200667 281869 200701 281897
rect 200729 281869 200763 281897
rect 200791 281869 200839 281897
rect 200529 281835 200839 281869
rect 200529 281807 200577 281835
rect 200605 281807 200639 281835
rect 200667 281807 200701 281835
rect 200729 281807 200763 281835
rect 200791 281807 200839 281835
rect 200529 281773 200839 281807
rect 200529 281745 200577 281773
rect 200605 281745 200639 281773
rect 200667 281745 200701 281773
rect 200729 281745 200763 281773
rect 200791 281745 200839 281773
rect 200529 272959 200839 281745
rect 200529 272931 200577 272959
rect 200605 272931 200639 272959
rect 200667 272931 200701 272959
rect 200729 272931 200763 272959
rect 200791 272931 200839 272959
rect 200529 272897 200839 272931
rect 200529 272869 200577 272897
rect 200605 272869 200639 272897
rect 200667 272869 200701 272897
rect 200729 272869 200763 272897
rect 200791 272869 200839 272897
rect 200529 272835 200839 272869
rect 200529 272807 200577 272835
rect 200605 272807 200639 272835
rect 200667 272807 200701 272835
rect 200729 272807 200763 272835
rect 200791 272807 200839 272835
rect 200529 272773 200839 272807
rect 200529 272745 200577 272773
rect 200605 272745 200639 272773
rect 200667 272745 200701 272773
rect 200729 272745 200763 272773
rect 200791 272745 200839 272773
rect 200529 263959 200839 272745
rect 200529 263931 200577 263959
rect 200605 263931 200639 263959
rect 200667 263931 200701 263959
rect 200729 263931 200763 263959
rect 200791 263931 200839 263959
rect 200529 263897 200839 263931
rect 200529 263869 200577 263897
rect 200605 263869 200639 263897
rect 200667 263869 200701 263897
rect 200729 263869 200763 263897
rect 200791 263869 200839 263897
rect 200529 263835 200839 263869
rect 200529 263807 200577 263835
rect 200605 263807 200639 263835
rect 200667 263807 200701 263835
rect 200729 263807 200763 263835
rect 200791 263807 200839 263835
rect 200529 263773 200839 263807
rect 200529 263745 200577 263773
rect 200605 263745 200639 263773
rect 200667 263745 200701 263773
rect 200729 263745 200763 263773
rect 200791 263745 200839 263773
rect 200529 254959 200839 263745
rect 200529 254931 200577 254959
rect 200605 254931 200639 254959
rect 200667 254931 200701 254959
rect 200729 254931 200763 254959
rect 200791 254931 200839 254959
rect 200529 254897 200839 254931
rect 200529 254869 200577 254897
rect 200605 254869 200639 254897
rect 200667 254869 200701 254897
rect 200729 254869 200763 254897
rect 200791 254869 200839 254897
rect 200529 254835 200839 254869
rect 200529 254807 200577 254835
rect 200605 254807 200639 254835
rect 200667 254807 200701 254835
rect 200729 254807 200763 254835
rect 200791 254807 200839 254835
rect 200529 254773 200839 254807
rect 200529 254745 200577 254773
rect 200605 254745 200639 254773
rect 200667 254745 200701 254773
rect 200729 254745 200763 254773
rect 200791 254745 200839 254773
rect 200529 254075 200839 254745
rect 202389 299670 202699 299718
rect 202389 299642 202437 299670
rect 202465 299642 202499 299670
rect 202527 299642 202561 299670
rect 202589 299642 202623 299670
rect 202651 299642 202699 299670
rect 202389 299608 202699 299642
rect 202389 299580 202437 299608
rect 202465 299580 202499 299608
rect 202527 299580 202561 299608
rect 202589 299580 202623 299608
rect 202651 299580 202699 299608
rect 202389 299546 202699 299580
rect 202389 299518 202437 299546
rect 202465 299518 202499 299546
rect 202527 299518 202561 299546
rect 202589 299518 202623 299546
rect 202651 299518 202699 299546
rect 202389 299484 202699 299518
rect 202389 299456 202437 299484
rect 202465 299456 202499 299484
rect 202527 299456 202561 299484
rect 202589 299456 202623 299484
rect 202651 299456 202699 299484
rect 202389 293959 202699 299456
rect 202389 293931 202437 293959
rect 202465 293931 202499 293959
rect 202527 293931 202561 293959
rect 202589 293931 202623 293959
rect 202651 293931 202699 293959
rect 202389 293897 202699 293931
rect 202389 293869 202437 293897
rect 202465 293869 202499 293897
rect 202527 293869 202561 293897
rect 202589 293869 202623 293897
rect 202651 293869 202699 293897
rect 202389 293835 202699 293869
rect 202389 293807 202437 293835
rect 202465 293807 202499 293835
rect 202527 293807 202561 293835
rect 202589 293807 202623 293835
rect 202651 293807 202699 293835
rect 202389 293773 202699 293807
rect 202389 293745 202437 293773
rect 202465 293745 202499 293773
rect 202527 293745 202561 293773
rect 202589 293745 202623 293773
rect 202651 293745 202699 293773
rect 202389 284959 202699 293745
rect 202389 284931 202437 284959
rect 202465 284931 202499 284959
rect 202527 284931 202561 284959
rect 202589 284931 202623 284959
rect 202651 284931 202699 284959
rect 202389 284897 202699 284931
rect 202389 284869 202437 284897
rect 202465 284869 202499 284897
rect 202527 284869 202561 284897
rect 202589 284869 202623 284897
rect 202651 284869 202699 284897
rect 202389 284835 202699 284869
rect 202389 284807 202437 284835
rect 202465 284807 202499 284835
rect 202527 284807 202561 284835
rect 202589 284807 202623 284835
rect 202651 284807 202699 284835
rect 202389 284773 202699 284807
rect 202389 284745 202437 284773
rect 202465 284745 202499 284773
rect 202527 284745 202561 284773
rect 202589 284745 202623 284773
rect 202651 284745 202699 284773
rect 202389 275959 202699 284745
rect 202389 275931 202437 275959
rect 202465 275931 202499 275959
rect 202527 275931 202561 275959
rect 202589 275931 202623 275959
rect 202651 275931 202699 275959
rect 202389 275897 202699 275931
rect 202389 275869 202437 275897
rect 202465 275869 202499 275897
rect 202527 275869 202561 275897
rect 202589 275869 202623 275897
rect 202651 275869 202699 275897
rect 202389 275835 202699 275869
rect 202389 275807 202437 275835
rect 202465 275807 202499 275835
rect 202527 275807 202561 275835
rect 202589 275807 202623 275835
rect 202651 275807 202699 275835
rect 202389 275773 202699 275807
rect 202389 275745 202437 275773
rect 202465 275745 202499 275773
rect 202527 275745 202561 275773
rect 202589 275745 202623 275773
rect 202651 275745 202699 275773
rect 202389 266959 202699 275745
rect 202389 266931 202437 266959
rect 202465 266931 202499 266959
rect 202527 266931 202561 266959
rect 202589 266931 202623 266959
rect 202651 266931 202699 266959
rect 202389 266897 202699 266931
rect 202389 266869 202437 266897
rect 202465 266869 202499 266897
rect 202527 266869 202561 266897
rect 202589 266869 202623 266897
rect 202651 266869 202699 266897
rect 202389 266835 202699 266869
rect 202389 266807 202437 266835
rect 202465 266807 202499 266835
rect 202527 266807 202561 266835
rect 202589 266807 202623 266835
rect 202651 266807 202699 266835
rect 202389 266773 202699 266807
rect 202389 266745 202437 266773
rect 202465 266745 202499 266773
rect 202527 266745 202561 266773
rect 202589 266745 202623 266773
rect 202651 266745 202699 266773
rect 202389 257959 202699 266745
rect 202389 257931 202437 257959
rect 202465 257931 202499 257959
rect 202527 257931 202561 257959
rect 202589 257931 202623 257959
rect 202651 257931 202699 257959
rect 202389 257897 202699 257931
rect 202389 257869 202437 257897
rect 202465 257869 202499 257897
rect 202527 257869 202561 257897
rect 202589 257869 202623 257897
rect 202651 257869 202699 257897
rect 202389 257835 202699 257869
rect 202389 257807 202437 257835
rect 202465 257807 202499 257835
rect 202527 257807 202561 257835
rect 202589 257807 202623 257835
rect 202651 257807 202699 257835
rect 202389 257773 202699 257807
rect 202389 257745 202437 257773
rect 202465 257745 202499 257773
rect 202527 257745 202561 257773
rect 202589 257745 202623 257773
rect 202651 257745 202699 257773
rect 202389 254075 202699 257745
rect 209529 299190 209839 299718
rect 209529 299162 209577 299190
rect 209605 299162 209639 299190
rect 209667 299162 209701 299190
rect 209729 299162 209763 299190
rect 209791 299162 209839 299190
rect 209529 299128 209839 299162
rect 209529 299100 209577 299128
rect 209605 299100 209639 299128
rect 209667 299100 209701 299128
rect 209729 299100 209763 299128
rect 209791 299100 209839 299128
rect 209529 299066 209839 299100
rect 209529 299038 209577 299066
rect 209605 299038 209639 299066
rect 209667 299038 209701 299066
rect 209729 299038 209763 299066
rect 209791 299038 209839 299066
rect 209529 299004 209839 299038
rect 209529 298976 209577 299004
rect 209605 298976 209639 299004
rect 209667 298976 209701 299004
rect 209729 298976 209763 299004
rect 209791 298976 209839 299004
rect 209529 290959 209839 298976
rect 209529 290931 209577 290959
rect 209605 290931 209639 290959
rect 209667 290931 209701 290959
rect 209729 290931 209763 290959
rect 209791 290931 209839 290959
rect 209529 290897 209839 290931
rect 209529 290869 209577 290897
rect 209605 290869 209639 290897
rect 209667 290869 209701 290897
rect 209729 290869 209763 290897
rect 209791 290869 209839 290897
rect 209529 290835 209839 290869
rect 209529 290807 209577 290835
rect 209605 290807 209639 290835
rect 209667 290807 209701 290835
rect 209729 290807 209763 290835
rect 209791 290807 209839 290835
rect 209529 290773 209839 290807
rect 209529 290745 209577 290773
rect 209605 290745 209639 290773
rect 209667 290745 209701 290773
rect 209729 290745 209763 290773
rect 209791 290745 209839 290773
rect 209529 281959 209839 290745
rect 209529 281931 209577 281959
rect 209605 281931 209639 281959
rect 209667 281931 209701 281959
rect 209729 281931 209763 281959
rect 209791 281931 209839 281959
rect 209529 281897 209839 281931
rect 209529 281869 209577 281897
rect 209605 281869 209639 281897
rect 209667 281869 209701 281897
rect 209729 281869 209763 281897
rect 209791 281869 209839 281897
rect 209529 281835 209839 281869
rect 209529 281807 209577 281835
rect 209605 281807 209639 281835
rect 209667 281807 209701 281835
rect 209729 281807 209763 281835
rect 209791 281807 209839 281835
rect 209529 281773 209839 281807
rect 209529 281745 209577 281773
rect 209605 281745 209639 281773
rect 209667 281745 209701 281773
rect 209729 281745 209763 281773
rect 209791 281745 209839 281773
rect 209529 272959 209839 281745
rect 209529 272931 209577 272959
rect 209605 272931 209639 272959
rect 209667 272931 209701 272959
rect 209729 272931 209763 272959
rect 209791 272931 209839 272959
rect 209529 272897 209839 272931
rect 209529 272869 209577 272897
rect 209605 272869 209639 272897
rect 209667 272869 209701 272897
rect 209729 272869 209763 272897
rect 209791 272869 209839 272897
rect 209529 272835 209839 272869
rect 209529 272807 209577 272835
rect 209605 272807 209639 272835
rect 209667 272807 209701 272835
rect 209729 272807 209763 272835
rect 209791 272807 209839 272835
rect 209529 272773 209839 272807
rect 209529 272745 209577 272773
rect 209605 272745 209639 272773
rect 209667 272745 209701 272773
rect 209729 272745 209763 272773
rect 209791 272745 209839 272773
rect 209529 263959 209839 272745
rect 209529 263931 209577 263959
rect 209605 263931 209639 263959
rect 209667 263931 209701 263959
rect 209729 263931 209763 263959
rect 209791 263931 209839 263959
rect 209529 263897 209839 263931
rect 209529 263869 209577 263897
rect 209605 263869 209639 263897
rect 209667 263869 209701 263897
rect 209729 263869 209763 263897
rect 209791 263869 209839 263897
rect 209529 263835 209839 263869
rect 209529 263807 209577 263835
rect 209605 263807 209639 263835
rect 209667 263807 209701 263835
rect 209729 263807 209763 263835
rect 209791 263807 209839 263835
rect 209529 263773 209839 263807
rect 209529 263745 209577 263773
rect 209605 263745 209639 263773
rect 209667 263745 209701 263773
rect 209729 263745 209763 263773
rect 209791 263745 209839 263773
rect 209529 254959 209839 263745
rect 209529 254931 209577 254959
rect 209605 254931 209639 254959
rect 209667 254931 209701 254959
rect 209729 254931 209763 254959
rect 209791 254931 209839 254959
rect 209529 254897 209839 254931
rect 209529 254869 209577 254897
rect 209605 254869 209639 254897
rect 209667 254869 209701 254897
rect 209729 254869 209763 254897
rect 209791 254869 209839 254897
rect 209529 254835 209839 254869
rect 209529 254807 209577 254835
rect 209605 254807 209639 254835
rect 209667 254807 209701 254835
rect 209729 254807 209763 254835
rect 209791 254807 209839 254835
rect 209529 254773 209839 254807
rect 209529 254745 209577 254773
rect 209605 254745 209639 254773
rect 209667 254745 209701 254773
rect 209729 254745 209763 254773
rect 209791 254745 209839 254773
rect 209529 254075 209839 254745
rect 211389 299670 211699 299718
rect 211389 299642 211437 299670
rect 211465 299642 211499 299670
rect 211527 299642 211561 299670
rect 211589 299642 211623 299670
rect 211651 299642 211699 299670
rect 211389 299608 211699 299642
rect 211389 299580 211437 299608
rect 211465 299580 211499 299608
rect 211527 299580 211561 299608
rect 211589 299580 211623 299608
rect 211651 299580 211699 299608
rect 211389 299546 211699 299580
rect 211389 299518 211437 299546
rect 211465 299518 211499 299546
rect 211527 299518 211561 299546
rect 211589 299518 211623 299546
rect 211651 299518 211699 299546
rect 211389 299484 211699 299518
rect 211389 299456 211437 299484
rect 211465 299456 211499 299484
rect 211527 299456 211561 299484
rect 211589 299456 211623 299484
rect 211651 299456 211699 299484
rect 211389 293959 211699 299456
rect 211389 293931 211437 293959
rect 211465 293931 211499 293959
rect 211527 293931 211561 293959
rect 211589 293931 211623 293959
rect 211651 293931 211699 293959
rect 211389 293897 211699 293931
rect 211389 293869 211437 293897
rect 211465 293869 211499 293897
rect 211527 293869 211561 293897
rect 211589 293869 211623 293897
rect 211651 293869 211699 293897
rect 211389 293835 211699 293869
rect 211389 293807 211437 293835
rect 211465 293807 211499 293835
rect 211527 293807 211561 293835
rect 211589 293807 211623 293835
rect 211651 293807 211699 293835
rect 211389 293773 211699 293807
rect 211389 293745 211437 293773
rect 211465 293745 211499 293773
rect 211527 293745 211561 293773
rect 211589 293745 211623 293773
rect 211651 293745 211699 293773
rect 211389 284959 211699 293745
rect 211389 284931 211437 284959
rect 211465 284931 211499 284959
rect 211527 284931 211561 284959
rect 211589 284931 211623 284959
rect 211651 284931 211699 284959
rect 211389 284897 211699 284931
rect 211389 284869 211437 284897
rect 211465 284869 211499 284897
rect 211527 284869 211561 284897
rect 211589 284869 211623 284897
rect 211651 284869 211699 284897
rect 211389 284835 211699 284869
rect 211389 284807 211437 284835
rect 211465 284807 211499 284835
rect 211527 284807 211561 284835
rect 211589 284807 211623 284835
rect 211651 284807 211699 284835
rect 211389 284773 211699 284807
rect 211389 284745 211437 284773
rect 211465 284745 211499 284773
rect 211527 284745 211561 284773
rect 211589 284745 211623 284773
rect 211651 284745 211699 284773
rect 211389 275959 211699 284745
rect 211389 275931 211437 275959
rect 211465 275931 211499 275959
rect 211527 275931 211561 275959
rect 211589 275931 211623 275959
rect 211651 275931 211699 275959
rect 211389 275897 211699 275931
rect 211389 275869 211437 275897
rect 211465 275869 211499 275897
rect 211527 275869 211561 275897
rect 211589 275869 211623 275897
rect 211651 275869 211699 275897
rect 211389 275835 211699 275869
rect 211389 275807 211437 275835
rect 211465 275807 211499 275835
rect 211527 275807 211561 275835
rect 211589 275807 211623 275835
rect 211651 275807 211699 275835
rect 211389 275773 211699 275807
rect 211389 275745 211437 275773
rect 211465 275745 211499 275773
rect 211527 275745 211561 275773
rect 211589 275745 211623 275773
rect 211651 275745 211699 275773
rect 211389 266959 211699 275745
rect 211389 266931 211437 266959
rect 211465 266931 211499 266959
rect 211527 266931 211561 266959
rect 211589 266931 211623 266959
rect 211651 266931 211699 266959
rect 211389 266897 211699 266931
rect 211389 266869 211437 266897
rect 211465 266869 211499 266897
rect 211527 266869 211561 266897
rect 211589 266869 211623 266897
rect 211651 266869 211699 266897
rect 211389 266835 211699 266869
rect 211389 266807 211437 266835
rect 211465 266807 211499 266835
rect 211527 266807 211561 266835
rect 211589 266807 211623 266835
rect 211651 266807 211699 266835
rect 211389 266773 211699 266807
rect 211389 266745 211437 266773
rect 211465 266745 211499 266773
rect 211527 266745 211561 266773
rect 211589 266745 211623 266773
rect 211651 266745 211699 266773
rect 211389 257959 211699 266745
rect 211389 257931 211437 257959
rect 211465 257931 211499 257959
rect 211527 257931 211561 257959
rect 211589 257931 211623 257959
rect 211651 257931 211699 257959
rect 211389 257897 211699 257931
rect 211389 257869 211437 257897
rect 211465 257869 211499 257897
rect 211527 257869 211561 257897
rect 211589 257869 211623 257897
rect 211651 257869 211699 257897
rect 211389 257835 211699 257869
rect 211389 257807 211437 257835
rect 211465 257807 211499 257835
rect 211527 257807 211561 257835
rect 211589 257807 211623 257835
rect 211651 257807 211699 257835
rect 211389 257773 211699 257807
rect 211389 257745 211437 257773
rect 211465 257745 211499 257773
rect 211527 257745 211561 257773
rect 211589 257745 211623 257773
rect 211651 257745 211699 257773
rect 211389 254075 211699 257745
rect 218529 299190 218839 299718
rect 218529 299162 218577 299190
rect 218605 299162 218639 299190
rect 218667 299162 218701 299190
rect 218729 299162 218763 299190
rect 218791 299162 218839 299190
rect 218529 299128 218839 299162
rect 218529 299100 218577 299128
rect 218605 299100 218639 299128
rect 218667 299100 218701 299128
rect 218729 299100 218763 299128
rect 218791 299100 218839 299128
rect 218529 299066 218839 299100
rect 218529 299038 218577 299066
rect 218605 299038 218639 299066
rect 218667 299038 218701 299066
rect 218729 299038 218763 299066
rect 218791 299038 218839 299066
rect 218529 299004 218839 299038
rect 218529 298976 218577 299004
rect 218605 298976 218639 299004
rect 218667 298976 218701 299004
rect 218729 298976 218763 299004
rect 218791 298976 218839 299004
rect 218529 290959 218839 298976
rect 218529 290931 218577 290959
rect 218605 290931 218639 290959
rect 218667 290931 218701 290959
rect 218729 290931 218763 290959
rect 218791 290931 218839 290959
rect 218529 290897 218839 290931
rect 218529 290869 218577 290897
rect 218605 290869 218639 290897
rect 218667 290869 218701 290897
rect 218729 290869 218763 290897
rect 218791 290869 218839 290897
rect 218529 290835 218839 290869
rect 218529 290807 218577 290835
rect 218605 290807 218639 290835
rect 218667 290807 218701 290835
rect 218729 290807 218763 290835
rect 218791 290807 218839 290835
rect 218529 290773 218839 290807
rect 218529 290745 218577 290773
rect 218605 290745 218639 290773
rect 218667 290745 218701 290773
rect 218729 290745 218763 290773
rect 218791 290745 218839 290773
rect 218529 281959 218839 290745
rect 218529 281931 218577 281959
rect 218605 281931 218639 281959
rect 218667 281931 218701 281959
rect 218729 281931 218763 281959
rect 218791 281931 218839 281959
rect 218529 281897 218839 281931
rect 218529 281869 218577 281897
rect 218605 281869 218639 281897
rect 218667 281869 218701 281897
rect 218729 281869 218763 281897
rect 218791 281869 218839 281897
rect 218529 281835 218839 281869
rect 218529 281807 218577 281835
rect 218605 281807 218639 281835
rect 218667 281807 218701 281835
rect 218729 281807 218763 281835
rect 218791 281807 218839 281835
rect 218529 281773 218839 281807
rect 218529 281745 218577 281773
rect 218605 281745 218639 281773
rect 218667 281745 218701 281773
rect 218729 281745 218763 281773
rect 218791 281745 218839 281773
rect 218529 272959 218839 281745
rect 218529 272931 218577 272959
rect 218605 272931 218639 272959
rect 218667 272931 218701 272959
rect 218729 272931 218763 272959
rect 218791 272931 218839 272959
rect 218529 272897 218839 272931
rect 218529 272869 218577 272897
rect 218605 272869 218639 272897
rect 218667 272869 218701 272897
rect 218729 272869 218763 272897
rect 218791 272869 218839 272897
rect 218529 272835 218839 272869
rect 218529 272807 218577 272835
rect 218605 272807 218639 272835
rect 218667 272807 218701 272835
rect 218729 272807 218763 272835
rect 218791 272807 218839 272835
rect 218529 272773 218839 272807
rect 218529 272745 218577 272773
rect 218605 272745 218639 272773
rect 218667 272745 218701 272773
rect 218729 272745 218763 272773
rect 218791 272745 218839 272773
rect 218529 263959 218839 272745
rect 218529 263931 218577 263959
rect 218605 263931 218639 263959
rect 218667 263931 218701 263959
rect 218729 263931 218763 263959
rect 218791 263931 218839 263959
rect 218529 263897 218839 263931
rect 218529 263869 218577 263897
rect 218605 263869 218639 263897
rect 218667 263869 218701 263897
rect 218729 263869 218763 263897
rect 218791 263869 218839 263897
rect 218529 263835 218839 263869
rect 218529 263807 218577 263835
rect 218605 263807 218639 263835
rect 218667 263807 218701 263835
rect 218729 263807 218763 263835
rect 218791 263807 218839 263835
rect 218529 263773 218839 263807
rect 218529 263745 218577 263773
rect 218605 263745 218639 263773
rect 218667 263745 218701 263773
rect 218729 263745 218763 263773
rect 218791 263745 218839 263773
rect 218529 254959 218839 263745
rect 218529 254931 218577 254959
rect 218605 254931 218639 254959
rect 218667 254931 218701 254959
rect 218729 254931 218763 254959
rect 218791 254931 218839 254959
rect 218529 254897 218839 254931
rect 218529 254869 218577 254897
rect 218605 254869 218639 254897
rect 218667 254869 218701 254897
rect 218729 254869 218763 254897
rect 218791 254869 218839 254897
rect 218529 254835 218839 254869
rect 218529 254807 218577 254835
rect 218605 254807 218639 254835
rect 218667 254807 218701 254835
rect 218729 254807 218763 254835
rect 218791 254807 218839 254835
rect 218529 254773 218839 254807
rect 218529 254745 218577 254773
rect 218605 254745 218639 254773
rect 218667 254745 218701 254773
rect 218729 254745 218763 254773
rect 218791 254745 218839 254773
rect 218529 254075 218839 254745
rect 220389 299670 220699 299718
rect 220389 299642 220437 299670
rect 220465 299642 220499 299670
rect 220527 299642 220561 299670
rect 220589 299642 220623 299670
rect 220651 299642 220699 299670
rect 220389 299608 220699 299642
rect 220389 299580 220437 299608
rect 220465 299580 220499 299608
rect 220527 299580 220561 299608
rect 220589 299580 220623 299608
rect 220651 299580 220699 299608
rect 220389 299546 220699 299580
rect 220389 299518 220437 299546
rect 220465 299518 220499 299546
rect 220527 299518 220561 299546
rect 220589 299518 220623 299546
rect 220651 299518 220699 299546
rect 220389 299484 220699 299518
rect 220389 299456 220437 299484
rect 220465 299456 220499 299484
rect 220527 299456 220561 299484
rect 220589 299456 220623 299484
rect 220651 299456 220699 299484
rect 220389 293959 220699 299456
rect 220389 293931 220437 293959
rect 220465 293931 220499 293959
rect 220527 293931 220561 293959
rect 220589 293931 220623 293959
rect 220651 293931 220699 293959
rect 220389 293897 220699 293931
rect 220389 293869 220437 293897
rect 220465 293869 220499 293897
rect 220527 293869 220561 293897
rect 220589 293869 220623 293897
rect 220651 293869 220699 293897
rect 220389 293835 220699 293869
rect 220389 293807 220437 293835
rect 220465 293807 220499 293835
rect 220527 293807 220561 293835
rect 220589 293807 220623 293835
rect 220651 293807 220699 293835
rect 220389 293773 220699 293807
rect 220389 293745 220437 293773
rect 220465 293745 220499 293773
rect 220527 293745 220561 293773
rect 220589 293745 220623 293773
rect 220651 293745 220699 293773
rect 220389 284959 220699 293745
rect 220389 284931 220437 284959
rect 220465 284931 220499 284959
rect 220527 284931 220561 284959
rect 220589 284931 220623 284959
rect 220651 284931 220699 284959
rect 220389 284897 220699 284931
rect 220389 284869 220437 284897
rect 220465 284869 220499 284897
rect 220527 284869 220561 284897
rect 220589 284869 220623 284897
rect 220651 284869 220699 284897
rect 220389 284835 220699 284869
rect 220389 284807 220437 284835
rect 220465 284807 220499 284835
rect 220527 284807 220561 284835
rect 220589 284807 220623 284835
rect 220651 284807 220699 284835
rect 220389 284773 220699 284807
rect 220389 284745 220437 284773
rect 220465 284745 220499 284773
rect 220527 284745 220561 284773
rect 220589 284745 220623 284773
rect 220651 284745 220699 284773
rect 220389 275959 220699 284745
rect 220389 275931 220437 275959
rect 220465 275931 220499 275959
rect 220527 275931 220561 275959
rect 220589 275931 220623 275959
rect 220651 275931 220699 275959
rect 220389 275897 220699 275931
rect 220389 275869 220437 275897
rect 220465 275869 220499 275897
rect 220527 275869 220561 275897
rect 220589 275869 220623 275897
rect 220651 275869 220699 275897
rect 220389 275835 220699 275869
rect 220389 275807 220437 275835
rect 220465 275807 220499 275835
rect 220527 275807 220561 275835
rect 220589 275807 220623 275835
rect 220651 275807 220699 275835
rect 220389 275773 220699 275807
rect 220389 275745 220437 275773
rect 220465 275745 220499 275773
rect 220527 275745 220561 275773
rect 220589 275745 220623 275773
rect 220651 275745 220699 275773
rect 220389 266959 220699 275745
rect 220389 266931 220437 266959
rect 220465 266931 220499 266959
rect 220527 266931 220561 266959
rect 220589 266931 220623 266959
rect 220651 266931 220699 266959
rect 220389 266897 220699 266931
rect 220389 266869 220437 266897
rect 220465 266869 220499 266897
rect 220527 266869 220561 266897
rect 220589 266869 220623 266897
rect 220651 266869 220699 266897
rect 220389 266835 220699 266869
rect 220389 266807 220437 266835
rect 220465 266807 220499 266835
rect 220527 266807 220561 266835
rect 220589 266807 220623 266835
rect 220651 266807 220699 266835
rect 220389 266773 220699 266807
rect 220389 266745 220437 266773
rect 220465 266745 220499 266773
rect 220527 266745 220561 266773
rect 220589 266745 220623 266773
rect 220651 266745 220699 266773
rect 220389 257959 220699 266745
rect 220389 257931 220437 257959
rect 220465 257931 220499 257959
rect 220527 257931 220561 257959
rect 220589 257931 220623 257959
rect 220651 257931 220699 257959
rect 220389 257897 220699 257931
rect 220389 257869 220437 257897
rect 220465 257869 220499 257897
rect 220527 257869 220561 257897
rect 220589 257869 220623 257897
rect 220651 257869 220699 257897
rect 220389 257835 220699 257869
rect 220389 257807 220437 257835
rect 220465 257807 220499 257835
rect 220527 257807 220561 257835
rect 220589 257807 220623 257835
rect 220651 257807 220699 257835
rect 220389 257773 220699 257807
rect 220389 257745 220437 257773
rect 220465 257745 220499 257773
rect 220527 257745 220561 257773
rect 220589 257745 220623 257773
rect 220651 257745 220699 257773
rect 220389 254075 220699 257745
rect 227529 299190 227839 299718
rect 227529 299162 227577 299190
rect 227605 299162 227639 299190
rect 227667 299162 227701 299190
rect 227729 299162 227763 299190
rect 227791 299162 227839 299190
rect 227529 299128 227839 299162
rect 227529 299100 227577 299128
rect 227605 299100 227639 299128
rect 227667 299100 227701 299128
rect 227729 299100 227763 299128
rect 227791 299100 227839 299128
rect 227529 299066 227839 299100
rect 227529 299038 227577 299066
rect 227605 299038 227639 299066
rect 227667 299038 227701 299066
rect 227729 299038 227763 299066
rect 227791 299038 227839 299066
rect 227529 299004 227839 299038
rect 227529 298976 227577 299004
rect 227605 298976 227639 299004
rect 227667 298976 227701 299004
rect 227729 298976 227763 299004
rect 227791 298976 227839 299004
rect 227529 290959 227839 298976
rect 227529 290931 227577 290959
rect 227605 290931 227639 290959
rect 227667 290931 227701 290959
rect 227729 290931 227763 290959
rect 227791 290931 227839 290959
rect 227529 290897 227839 290931
rect 227529 290869 227577 290897
rect 227605 290869 227639 290897
rect 227667 290869 227701 290897
rect 227729 290869 227763 290897
rect 227791 290869 227839 290897
rect 227529 290835 227839 290869
rect 227529 290807 227577 290835
rect 227605 290807 227639 290835
rect 227667 290807 227701 290835
rect 227729 290807 227763 290835
rect 227791 290807 227839 290835
rect 227529 290773 227839 290807
rect 227529 290745 227577 290773
rect 227605 290745 227639 290773
rect 227667 290745 227701 290773
rect 227729 290745 227763 290773
rect 227791 290745 227839 290773
rect 227529 281959 227839 290745
rect 227529 281931 227577 281959
rect 227605 281931 227639 281959
rect 227667 281931 227701 281959
rect 227729 281931 227763 281959
rect 227791 281931 227839 281959
rect 227529 281897 227839 281931
rect 227529 281869 227577 281897
rect 227605 281869 227639 281897
rect 227667 281869 227701 281897
rect 227729 281869 227763 281897
rect 227791 281869 227839 281897
rect 227529 281835 227839 281869
rect 227529 281807 227577 281835
rect 227605 281807 227639 281835
rect 227667 281807 227701 281835
rect 227729 281807 227763 281835
rect 227791 281807 227839 281835
rect 227529 281773 227839 281807
rect 227529 281745 227577 281773
rect 227605 281745 227639 281773
rect 227667 281745 227701 281773
rect 227729 281745 227763 281773
rect 227791 281745 227839 281773
rect 227529 272959 227839 281745
rect 227529 272931 227577 272959
rect 227605 272931 227639 272959
rect 227667 272931 227701 272959
rect 227729 272931 227763 272959
rect 227791 272931 227839 272959
rect 227529 272897 227839 272931
rect 227529 272869 227577 272897
rect 227605 272869 227639 272897
rect 227667 272869 227701 272897
rect 227729 272869 227763 272897
rect 227791 272869 227839 272897
rect 227529 272835 227839 272869
rect 227529 272807 227577 272835
rect 227605 272807 227639 272835
rect 227667 272807 227701 272835
rect 227729 272807 227763 272835
rect 227791 272807 227839 272835
rect 227529 272773 227839 272807
rect 227529 272745 227577 272773
rect 227605 272745 227639 272773
rect 227667 272745 227701 272773
rect 227729 272745 227763 272773
rect 227791 272745 227839 272773
rect 227529 263959 227839 272745
rect 227529 263931 227577 263959
rect 227605 263931 227639 263959
rect 227667 263931 227701 263959
rect 227729 263931 227763 263959
rect 227791 263931 227839 263959
rect 227529 263897 227839 263931
rect 227529 263869 227577 263897
rect 227605 263869 227639 263897
rect 227667 263869 227701 263897
rect 227729 263869 227763 263897
rect 227791 263869 227839 263897
rect 227529 263835 227839 263869
rect 227529 263807 227577 263835
rect 227605 263807 227639 263835
rect 227667 263807 227701 263835
rect 227729 263807 227763 263835
rect 227791 263807 227839 263835
rect 227529 263773 227839 263807
rect 227529 263745 227577 263773
rect 227605 263745 227639 263773
rect 227667 263745 227701 263773
rect 227729 263745 227763 263773
rect 227791 263745 227839 263773
rect 227529 254959 227839 263745
rect 227529 254931 227577 254959
rect 227605 254931 227639 254959
rect 227667 254931 227701 254959
rect 227729 254931 227763 254959
rect 227791 254931 227839 254959
rect 227529 254897 227839 254931
rect 227529 254869 227577 254897
rect 227605 254869 227639 254897
rect 227667 254869 227701 254897
rect 227729 254869 227763 254897
rect 227791 254869 227839 254897
rect 227529 254835 227839 254869
rect 227529 254807 227577 254835
rect 227605 254807 227639 254835
rect 227667 254807 227701 254835
rect 227729 254807 227763 254835
rect 227791 254807 227839 254835
rect 227529 254773 227839 254807
rect 227529 254745 227577 254773
rect 227605 254745 227639 254773
rect 227667 254745 227701 254773
rect 227729 254745 227763 254773
rect 227791 254745 227839 254773
rect 227529 254075 227839 254745
rect 229389 299670 229699 299718
rect 229389 299642 229437 299670
rect 229465 299642 229499 299670
rect 229527 299642 229561 299670
rect 229589 299642 229623 299670
rect 229651 299642 229699 299670
rect 229389 299608 229699 299642
rect 229389 299580 229437 299608
rect 229465 299580 229499 299608
rect 229527 299580 229561 299608
rect 229589 299580 229623 299608
rect 229651 299580 229699 299608
rect 229389 299546 229699 299580
rect 229389 299518 229437 299546
rect 229465 299518 229499 299546
rect 229527 299518 229561 299546
rect 229589 299518 229623 299546
rect 229651 299518 229699 299546
rect 229389 299484 229699 299518
rect 229389 299456 229437 299484
rect 229465 299456 229499 299484
rect 229527 299456 229561 299484
rect 229589 299456 229623 299484
rect 229651 299456 229699 299484
rect 229389 293959 229699 299456
rect 229389 293931 229437 293959
rect 229465 293931 229499 293959
rect 229527 293931 229561 293959
rect 229589 293931 229623 293959
rect 229651 293931 229699 293959
rect 229389 293897 229699 293931
rect 229389 293869 229437 293897
rect 229465 293869 229499 293897
rect 229527 293869 229561 293897
rect 229589 293869 229623 293897
rect 229651 293869 229699 293897
rect 229389 293835 229699 293869
rect 229389 293807 229437 293835
rect 229465 293807 229499 293835
rect 229527 293807 229561 293835
rect 229589 293807 229623 293835
rect 229651 293807 229699 293835
rect 229389 293773 229699 293807
rect 229389 293745 229437 293773
rect 229465 293745 229499 293773
rect 229527 293745 229561 293773
rect 229589 293745 229623 293773
rect 229651 293745 229699 293773
rect 229389 284959 229699 293745
rect 229389 284931 229437 284959
rect 229465 284931 229499 284959
rect 229527 284931 229561 284959
rect 229589 284931 229623 284959
rect 229651 284931 229699 284959
rect 229389 284897 229699 284931
rect 229389 284869 229437 284897
rect 229465 284869 229499 284897
rect 229527 284869 229561 284897
rect 229589 284869 229623 284897
rect 229651 284869 229699 284897
rect 229389 284835 229699 284869
rect 229389 284807 229437 284835
rect 229465 284807 229499 284835
rect 229527 284807 229561 284835
rect 229589 284807 229623 284835
rect 229651 284807 229699 284835
rect 229389 284773 229699 284807
rect 229389 284745 229437 284773
rect 229465 284745 229499 284773
rect 229527 284745 229561 284773
rect 229589 284745 229623 284773
rect 229651 284745 229699 284773
rect 229389 275959 229699 284745
rect 229389 275931 229437 275959
rect 229465 275931 229499 275959
rect 229527 275931 229561 275959
rect 229589 275931 229623 275959
rect 229651 275931 229699 275959
rect 229389 275897 229699 275931
rect 229389 275869 229437 275897
rect 229465 275869 229499 275897
rect 229527 275869 229561 275897
rect 229589 275869 229623 275897
rect 229651 275869 229699 275897
rect 229389 275835 229699 275869
rect 229389 275807 229437 275835
rect 229465 275807 229499 275835
rect 229527 275807 229561 275835
rect 229589 275807 229623 275835
rect 229651 275807 229699 275835
rect 229389 275773 229699 275807
rect 229389 275745 229437 275773
rect 229465 275745 229499 275773
rect 229527 275745 229561 275773
rect 229589 275745 229623 275773
rect 229651 275745 229699 275773
rect 229389 266959 229699 275745
rect 229389 266931 229437 266959
rect 229465 266931 229499 266959
rect 229527 266931 229561 266959
rect 229589 266931 229623 266959
rect 229651 266931 229699 266959
rect 229389 266897 229699 266931
rect 229389 266869 229437 266897
rect 229465 266869 229499 266897
rect 229527 266869 229561 266897
rect 229589 266869 229623 266897
rect 229651 266869 229699 266897
rect 229389 266835 229699 266869
rect 229389 266807 229437 266835
rect 229465 266807 229499 266835
rect 229527 266807 229561 266835
rect 229589 266807 229623 266835
rect 229651 266807 229699 266835
rect 229389 266773 229699 266807
rect 229389 266745 229437 266773
rect 229465 266745 229499 266773
rect 229527 266745 229561 266773
rect 229589 266745 229623 266773
rect 229651 266745 229699 266773
rect 229389 257959 229699 266745
rect 229389 257931 229437 257959
rect 229465 257931 229499 257959
rect 229527 257931 229561 257959
rect 229589 257931 229623 257959
rect 229651 257931 229699 257959
rect 229389 257897 229699 257931
rect 229389 257869 229437 257897
rect 229465 257869 229499 257897
rect 229527 257869 229561 257897
rect 229589 257869 229623 257897
rect 229651 257869 229699 257897
rect 229389 257835 229699 257869
rect 229389 257807 229437 257835
rect 229465 257807 229499 257835
rect 229527 257807 229561 257835
rect 229589 257807 229623 257835
rect 229651 257807 229699 257835
rect 229389 257773 229699 257807
rect 229389 257745 229437 257773
rect 229465 257745 229499 257773
rect 229527 257745 229561 257773
rect 229589 257745 229623 257773
rect 229651 257745 229699 257773
rect 229389 254075 229699 257745
rect 236529 299190 236839 299718
rect 236529 299162 236577 299190
rect 236605 299162 236639 299190
rect 236667 299162 236701 299190
rect 236729 299162 236763 299190
rect 236791 299162 236839 299190
rect 236529 299128 236839 299162
rect 236529 299100 236577 299128
rect 236605 299100 236639 299128
rect 236667 299100 236701 299128
rect 236729 299100 236763 299128
rect 236791 299100 236839 299128
rect 236529 299066 236839 299100
rect 236529 299038 236577 299066
rect 236605 299038 236639 299066
rect 236667 299038 236701 299066
rect 236729 299038 236763 299066
rect 236791 299038 236839 299066
rect 236529 299004 236839 299038
rect 236529 298976 236577 299004
rect 236605 298976 236639 299004
rect 236667 298976 236701 299004
rect 236729 298976 236763 299004
rect 236791 298976 236839 299004
rect 236529 290959 236839 298976
rect 236529 290931 236577 290959
rect 236605 290931 236639 290959
rect 236667 290931 236701 290959
rect 236729 290931 236763 290959
rect 236791 290931 236839 290959
rect 236529 290897 236839 290931
rect 236529 290869 236577 290897
rect 236605 290869 236639 290897
rect 236667 290869 236701 290897
rect 236729 290869 236763 290897
rect 236791 290869 236839 290897
rect 236529 290835 236839 290869
rect 236529 290807 236577 290835
rect 236605 290807 236639 290835
rect 236667 290807 236701 290835
rect 236729 290807 236763 290835
rect 236791 290807 236839 290835
rect 236529 290773 236839 290807
rect 236529 290745 236577 290773
rect 236605 290745 236639 290773
rect 236667 290745 236701 290773
rect 236729 290745 236763 290773
rect 236791 290745 236839 290773
rect 236529 281959 236839 290745
rect 236529 281931 236577 281959
rect 236605 281931 236639 281959
rect 236667 281931 236701 281959
rect 236729 281931 236763 281959
rect 236791 281931 236839 281959
rect 236529 281897 236839 281931
rect 236529 281869 236577 281897
rect 236605 281869 236639 281897
rect 236667 281869 236701 281897
rect 236729 281869 236763 281897
rect 236791 281869 236839 281897
rect 236529 281835 236839 281869
rect 236529 281807 236577 281835
rect 236605 281807 236639 281835
rect 236667 281807 236701 281835
rect 236729 281807 236763 281835
rect 236791 281807 236839 281835
rect 236529 281773 236839 281807
rect 236529 281745 236577 281773
rect 236605 281745 236639 281773
rect 236667 281745 236701 281773
rect 236729 281745 236763 281773
rect 236791 281745 236839 281773
rect 236529 272959 236839 281745
rect 236529 272931 236577 272959
rect 236605 272931 236639 272959
rect 236667 272931 236701 272959
rect 236729 272931 236763 272959
rect 236791 272931 236839 272959
rect 236529 272897 236839 272931
rect 236529 272869 236577 272897
rect 236605 272869 236639 272897
rect 236667 272869 236701 272897
rect 236729 272869 236763 272897
rect 236791 272869 236839 272897
rect 236529 272835 236839 272869
rect 236529 272807 236577 272835
rect 236605 272807 236639 272835
rect 236667 272807 236701 272835
rect 236729 272807 236763 272835
rect 236791 272807 236839 272835
rect 236529 272773 236839 272807
rect 236529 272745 236577 272773
rect 236605 272745 236639 272773
rect 236667 272745 236701 272773
rect 236729 272745 236763 272773
rect 236791 272745 236839 272773
rect 236529 263959 236839 272745
rect 236529 263931 236577 263959
rect 236605 263931 236639 263959
rect 236667 263931 236701 263959
rect 236729 263931 236763 263959
rect 236791 263931 236839 263959
rect 236529 263897 236839 263931
rect 236529 263869 236577 263897
rect 236605 263869 236639 263897
rect 236667 263869 236701 263897
rect 236729 263869 236763 263897
rect 236791 263869 236839 263897
rect 236529 263835 236839 263869
rect 236529 263807 236577 263835
rect 236605 263807 236639 263835
rect 236667 263807 236701 263835
rect 236729 263807 236763 263835
rect 236791 263807 236839 263835
rect 236529 263773 236839 263807
rect 236529 263745 236577 263773
rect 236605 263745 236639 263773
rect 236667 263745 236701 263773
rect 236729 263745 236763 263773
rect 236791 263745 236839 263773
rect 236529 254959 236839 263745
rect 236529 254931 236577 254959
rect 236605 254931 236639 254959
rect 236667 254931 236701 254959
rect 236729 254931 236763 254959
rect 236791 254931 236839 254959
rect 236529 254897 236839 254931
rect 236529 254869 236577 254897
rect 236605 254869 236639 254897
rect 236667 254869 236701 254897
rect 236729 254869 236763 254897
rect 236791 254869 236839 254897
rect 236529 254835 236839 254869
rect 236529 254807 236577 254835
rect 236605 254807 236639 254835
rect 236667 254807 236701 254835
rect 236729 254807 236763 254835
rect 236791 254807 236839 254835
rect 236529 254773 236839 254807
rect 236529 254745 236577 254773
rect 236605 254745 236639 254773
rect 236667 254745 236701 254773
rect 236729 254745 236763 254773
rect 236791 254745 236839 254773
rect 236529 254075 236839 254745
rect 238389 299670 238699 299718
rect 238389 299642 238437 299670
rect 238465 299642 238499 299670
rect 238527 299642 238561 299670
rect 238589 299642 238623 299670
rect 238651 299642 238699 299670
rect 238389 299608 238699 299642
rect 238389 299580 238437 299608
rect 238465 299580 238499 299608
rect 238527 299580 238561 299608
rect 238589 299580 238623 299608
rect 238651 299580 238699 299608
rect 238389 299546 238699 299580
rect 238389 299518 238437 299546
rect 238465 299518 238499 299546
rect 238527 299518 238561 299546
rect 238589 299518 238623 299546
rect 238651 299518 238699 299546
rect 238389 299484 238699 299518
rect 238389 299456 238437 299484
rect 238465 299456 238499 299484
rect 238527 299456 238561 299484
rect 238589 299456 238623 299484
rect 238651 299456 238699 299484
rect 238389 293959 238699 299456
rect 238389 293931 238437 293959
rect 238465 293931 238499 293959
rect 238527 293931 238561 293959
rect 238589 293931 238623 293959
rect 238651 293931 238699 293959
rect 238389 293897 238699 293931
rect 238389 293869 238437 293897
rect 238465 293869 238499 293897
rect 238527 293869 238561 293897
rect 238589 293869 238623 293897
rect 238651 293869 238699 293897
rect 238389 293835 238699 293869
rect 238389 293807 238437 293835
rect 238465 293807 238499 293835
rect 238527 293807 238561 293835
rect 238589 293807 238623 293835
rect 238651 293807 238699 293835
rect 238389 293773 238699 293807
rect 238389 293745 238437 293773
rect 238465 293745 238499 293773
rect 238527 293745 238561 293773
rect 238589 293745 238623 293773
rect 238651 293745 238699 293773
rect 238389 284959 238699 293745
rect 238389 284931 238437 284959
rect 238465 284931 238499 284959
rect 238527 284931 238561 284959
rect 238589 284931 238623 284959
rect 238651 284931 238699 284959
rect 238389 284897 238699 284931
rect 238389 284869 238437 284897
rect 238465 284869 238499 284897
rect 238527 284869 238561 284897
rect 238589 284869 238623 284897
rect 238651 284869 238699 284897
rect 238389 284835 238699 284869
rect 238389 284807 238437 284835
rect 238465 284807 238499 284835
rect 238527 284807 238561 284835
rect 238589 284807 238623 284835
rect 238651 284807 238699 284835
rect 238389 284773 238699 284807
rect 238389 284745 238437 284773
rect 238465 284745 238499 284773
rect 238527 284745 238561 284773
rect 238589 284745 238623 284773
rect 238651 284745 238699 284773
rect 238389 275959 238699 284745
rect 238389 275931 238437 275959
rect 238465 275931 238499 275959
rect 238527 275931 238561 275959
rect 238589 275931 238623 275959
rect 238651 275931 238699 275959
rect 238389 275897 238699 275931
rect 238389 275869 238437 275897
rect 238465 275869 238499 275897
rect 238527 275869 238561 275897
rect 238589 275869 238623 275897
rect 238651 275869 238699 275897
rect 238389 275835 238699 275869
rect 238389 275807 238437 275835
rect 238465 275807 238499 275835
rect 238527 275807 238561 275835
rect 238589 275807 238623 275835
rect 238651 275807 238699 275835
rect 238389 275773 238699 275807
rect 238389 275745 238437 275773
rect 238465 275745 238499 275773
rect 238527 275745 238561 275773
rect 238589 275745 238623 275773
rect 238651 275745 238699 275773
rect 238389 266959 238699 275745
rect 238389 266931 238437 266959
rect 238465 266931 238499 266959
rect 238527 266931 238561 266959
rect 238589 266931 238623 266959
rect 238651 266931 238699 266959
rect 238389 266897 238699 266931
rect 238389 266869 238437 266897
rect 238465 266869 238499 266897
rect 238527 266869 238561 266897
rect 238589 266869 238623 266897
rect 238651 266869 238699 266897
rect 238389 266835 238699 266869
rect 238389 266807 238437 266835
rect 238465 266807 238499 266835
rect 238527 266807 238561 266835
rect 238589 266807 238623 266835
rect 238651 266807 238699 266835
rect 238389 266773 238699 266807
rect 238389 266745 238437 266773
rect 238465 266745 238499 266773
rect 238527 266745 238561 266773
rect 238589 266745 238623 266773
rect 238651 266745 238699 266773
rect 238389 257959 238699 266745
rect 238389 257931 238437 257959
rect 238465 257931 238499 257959
rect 238527 257931 238561 257959
rect 238589 257931 238623 257959
rect 238651 257931 238699 257959
rect 238389 257897 238699 257931
rect 238389 257869 238437 257897
rect 238465 257869 238499 257897
rect 238527 257869 238561 257897
rect 238589 257869 238623 257897
rect 238651 257869 238699 257897
rect 238389 257835 238699 257869
rect 238389 257807 238437 257835
rect 238465 257807 238499 257835
rect 238527 257807 238561 257835
rect 238589 257807 238623 257835
rect 238651 257807 238699 257835
rect 238389 257773 238699 257807
rect 238389 257745 238437 257773
rect 238465 257745 238499 257773
rect 238527 257745 238561 257773
rect 238589 257745 238623 257773
rect 238651 257745 238699 257773
rect 238389 254075 238699 257745
rect 245529 299190 245839 299718
rect 245529 299162 245577 299190
rect 245605 299162 245639 299190
rect 245667 299162 245701 299190
rect 245729 299162 245763 299190
rect 245791 299162 245839 299190
rect 245529 299128 245839 299162
rect 245529 299100 245577 299128
rect 245605 299100 245639 299128
rect 245667 299100 245701 299128
rect 245729 299100 245763 299128
rect 245791 299100 245839 299128
rect 245529 299066 245839 299100
rect 245529 299038 245577 299066
rect 245605 299038 245639 299066
rect 245667 299038 245701 299066
rect 245729 299038 245763 299066
rect 245791 299038 245839 299066
rect 245529 299004 245839 299038
rect 245529 298976 245577 299004
rect 245605 298976 245639 299004
rect 245667 298976 245701 299004
rect 245729 298976 245763 299004
rect 245791 298976 245839 299004
rect 245529 290959 245839 298976
rect 245529 290931 245577 290959
rect 245605 290931 245639 290959
rect 245667 290931 245701 290959
rect 245729 290931 245763 290959
rect 245791 290931 245839 290959
rect 245529 290897 245839 290931
rect 245529 290869 245577 290897
rect 245605 290869 245639 290897
rect 245667 290869 245701 290897
rect 245729 290869 245763 290897
rect 245791 290869 245839 290897
rect 245529 290835 245839 290869
rect 245529 290807 245577 290835
rect 245605 290807 245639 290835
rect 245667 290807 245701 290835
rect 245729 290807 245763 290835
rect 245791 290807 245839 290835
rect 245529 290773 245839 290807
rect 245529 290745 245577 290773
rect 245605 290745 245639 290773
rect 245667 290745 245701 290773
rect 245729 290745 245763 290773
rect 245791 290745 245839 290773
rect 245529 281959 245839 290745
rect 245529 281931 245577 281959
rect 245605 281931 245639 281959
rect 245667 281931 245701 281959
rect 245729 281931 245763 281959
rect 245791 281931 245839 281959
rect 245529 281897 245839 281931
rect 245529 281869 245577 281897
rect 245605 281869 245639 281897
rect 245667 281869 245701 281897
rect 245729 281869 245763 281897
rect 245791 281869 245839 281897
rect 245529 281835 245839 281869
rect 245529 281807 245577 281835
rect 245605 281807 245639 281835
rect 245667 281807 245701 281835
rect 245729 281807 245763 281835
rect 245791 281807 245839 281835
rect 245529 281773 245839 281807
rect 245529 281745 245577 281773
rect 245605 281745 245639 281773
rect 245667 281745 245701 281773
rect 245729 281745 245763 281773
rect 245791 281745 245839 281773
rect 245529 272959 245839 281745
rect 245529 272931 245577 272959
rect 245605 272931 245639 272959
rect 245667 272931 245701 272959
rect 245729 272931 245763 272959
rect 245791 272931 245839 272959
rect 245529 272897 245839 272931
rect 245529 272869 245577 272897
rect 245605 272869 245639 272897
rect 245667 272869 245701 272897
rect 245729 272869 245763 272897
rect 245791 272869 245839 272897
rect 245529 272835 245839 272869
rect 245529 272807 245577 272835
rect 245605 272807 245639 272835
rect 245667 272807 245701 272835
rect 245729 272807 245763 272835
rect 245791 272807 245839 272835
rect 245529 272773 245839 272807
rect 245529 272745 245577 272773
rect 245605 272745 245639 272773
rect 245667 272745 245701 272773
rect 245729 272745 245763 272773
rect 245791 272745 245839 272773
rect 245529 263959 245839 272745
rect 245529 263931 245577 263959
rect 245605 263931 245639 263959
rect 245667 263931 245701 263959
rect 245729 263931 245763 263959
rect 245791 263931 245839 263959
rect 245529 263897 245839 263931
rect 245529 263869 245577 263897
rect 245605 263869 245639 263897
rect 245667 263869 245701 263897
rect 245729 263869 245763 263897
rect 245791 263869 245839 263897
rect 245529 263835 245839 263869
rect 245529 263807 245577 263835
rect 245605 263807 245639 263835
rect 245667 263807 245701 263835
rect 245729 263807 245763 263835
rect 245791 263807 245839 263835
rect 245529 263773 245839 263807
rect 245529 263745 245577 263773
rect 245605 263745 245639 263773
rect 245667 263745 245701 263773
rect 245729 263745 245763 263773
rect 245791 263745 245839 263773
rect 245529 254959 245839 263745
rect 245529 254931 245577 254959
rect 245605 254931 245639 254959
rect 245667 254931 245701 254959
rect 245729 254931 245763 254959
rect 245791 254931 245839 254959
rect 245529 254897 245839 254931
rect 245529 254869 245577 254897
rect 245605 254869 245639 254897
rect 245667 254869 245701 254897
rect 245729 254869 245763 254897
rect 245791 254869 245839 254897
rect 245529 254835 245839 254869
rect 245529 254807 245577 254835
rect 245605 254807 245639 254835
rect 245667 254807 245701 254835
rect 245729 254807 245763 254835
rect 245791 254807 245839 254835
rect 245529 254773 245839 254807
rect 245529 254745 245577 254773
rect 245605 254745 245639 254773
rect 245667 254745 245701 254773
rect 245729 254745 245763 254773
rect 245791 254745 245839 254773
rect 245529 254075 245839 254745
rect 247389 299670 247699 299718
rect 247389 299642 247437 299670
rect 247465 299642 247499 299670
rect 247527 299642 247561 299670
rect 247589 299642 247623 299670
rect 247651 299642 247699 299670
rect 247389 299608 247699 299642
rect 247389 299580 247437 299608
rect 247465 299580 247499 299608
rect 247527 299580 247561 299608
rect 247589 299580 247623 299608
rect 247651 299580 247699 299608
rect 247389 299546 247699 299580
rect 247389 299518 247437 299546
rect 247465 299518 247499 299546
rect 247527 299518 247561 299546
rect 247589 299518 247623 299546
rect 247651 299518 247699 299546
rect 247389 299484 247699 299518
rect 247389 299456 247437 299484
rect 247465 299456 247499 299484
rect 247527 299456 247561 299484
rect 247589 299456 247623 299484
rect 247651 299456 247699 299484
rect 247389 293959 247699 299456
rect 247389 293931 247437 293959
rect 247465 293931 247499 293959
rect 247527 293931 247561 293959
rect 247589 293931 247623 293959
rect 247651 293931 247699 293959
rect 247389 293897 247699 293931
rect 247389 293869 247437 293897
rect 247465 293869 247499 293897
rect 247527 293869 247561 293897
rect 247589 293869 247623 293897
rect 247651 293869 247699 293897
rect 247389 293835 247699 293869
rect 247389 293807 247437 293835
rect 247465 293807 247499 293835
rect 247527 293807 247561 293835
rect 247589 293807 247623 293835
rect 247651 293807 247699 293835
rect 247389 293773 247699 293807
rect 247389 293745 247437 293773
rect 247465 293745 247499 293773
rect 247527 293745 247561 293773
rect 247589 293745 247623 293773
rect 247651 293745 247699 293773
rect 247389 284959 247699 293745
rect 247389 284931 247437 284959
rect 247465 284931 247499 284959
rect 247527 284931 247561 284959
rect 247589 284931 247623 284959
rect 247651 284931 247699 284959
rect 247389 284897 247699 284931
rect 247389 284869 247437 284897
rect 247465 284869 247499 284897
rect 247527 284869 247561 284897
rect 247589 284869 247623 284897
rect 247651 284869 247699 284897
rect 247389 284835 247699 284869
rect 247389 284807 247437 284835
rect 247465 284807 247499 284835
rect 247527 284807 247561 284835
rect 247589 284807 247623 284835
rect 247651 284807 247699 284835
rect 247389 284773 247699 284807
rect 247389 284745 247437 284773
rect 247465 284745 247499 284773
rect 247527 284745 247561 284773
rect 247589 284745 247623 284773
rect 247651 284745 247699 284773
rect 247389 275959 247699 284745
rect 247389 275931 247437 275959
rect 247465 275931 247499 275959
rect 247527 275931 247561 275959
rect 247589 275931 247623 275959
rect 247651 275931 247699 275959
rect 247389 275897 247699 275931
rect 247389 275869 247437 275897
rect 247465 275869 247499 275897
rect 247527 275869 247561 275897
rect 247589 275869 247623 275897
rect 247651 275869 247699 275897
rect 247389 275835 247699 275869
rect 247389 275807 247437 275835
rect 247465 275807 247499 275835
rect 247527 275807 247561 275835
rect 247589 275807 247623 275835
rect 247651 275807 247699 275835
rect 247389 275773 247699 275807
rect 247389 275745 247437 275773
rect 247465 275745 247499 275773
rect 247527 275745 247561 275773
rect 247589 275745 247623 275773
rect 247651 275745 247699 275773
rect 247389 266959 247699 275745
rect 247389 266931 247437 266959
rect 247465 266931 247499 266959
rect 247527 266931 247561 266959
rect 247589 266931 247623 266959
rect 247651 266931 247699 266959
rect 247389 266897 247699 266931
rect 247389 266869 247437 266897
rect 247465 266869 247499 266897
rect 247527 266869 247561 266897
rect 247589 266869 247623 266897
rect 247651 266869 247699 266897
rect 247389 266835 247699 266869
rect 247389 266807 247437 266835
rect 247465 266807 247499 266835
rect 247527 266807 247561 266835
rect 247589 266807 247623 266835
rect 247651 266807 247699 266835
rect 247389 266773 247699 266807
rect 247389 266745 247437 266773
rect 247465 266745 247499 266773
rect 247527 266745 247561 266773
rect 247589 266745 247623 266773
rect 247651 266745 247699 266773
rect 247389 257959 247699 266745
rect 247389 257931 247437 257959
rect 247465 257931 247499 257959
rect 247527 257931 247561 257959
rect 247589 257931 247623 257959
rect 247651 257931 247699 257959
rect 247389 257897 247699 257931
rect 247389 257869 247437 257897
rect 247465 257869 247499 257897
rect 247527 257869 247561 257897
rect 247589 257869 247623 257897
rect 247651 257869 247699 257897
rect 247389 257835 247699 257869
rect 247389 257807 247437 257835
rect 247465 257807 247499 257835
rect 247527 257807 247561 257835
rect 247589 257807 247623 257835
rect 247651 257807 247699 257835
rect 247389 257773 247699 257807
rect 247389 257745 247437 257773
rect 247465 257745 247499 257773
rect 247527 257745 247561 257773
rect 247589 257745 247623 257773
rect 247651 257745 247699 257773
rect 247389 254394 247699 257745
rect 254529 299190 254839 299718
rect 254529 299162 254577 299190
rect 254605 299162 254639 299190
rect 254667 299162 254701 299190
rect 254729 299162 254763 299190
rect 254791 299162 254839 299190
rect 254529 299128 254839 299162
rect 254529 299100 254577 299128
rect 254605 299100 254639 299128
rect 254667 299100 254701 299128
rect 254729 299100 254763 299128
rect 254791 299100 254839 299128
rect 254529 299066 254839 299100
rect 254529 299038 254577 299066
rect 254605 299038 254639 299066
rect 254667 299038 254701 299066
rect 254729 299038 254763 299066
rect 254791 299038 254839 299066
rect 254529 299004 254839 299038
rect 254529 298976 254577 299004
rect 254605 298976 254639 299004
rect 254667 298976 254701 299004
rect 254729 298976 254763 299004
rect 254791 298976 254839 299004
rect 254529 290959 254839 298976
rect 254529 290931 254577 290959
rect 254605 290931 254639 290959
rect 254667 290931 254701 290959
rect 254729 290931 254763 290959
rect 254791 290931 254839 290959
rect 254529 290897 254839 290931
rect 254529 290869 254577 290897
rect 254605 290869 254639 290897
rect 254667 290869 254701 290897
rect 254729 290869 254763 290897
rect 254791 290869 254839 290897
rect 254529 290835 254839 290869
rect 254529 290807 254577 290835
rect 254605 290807 254639 290835
rect 254667 290807 254701 290835
rect 254729 290807 254763 290835
rect 254791 290807 254839 290835
rect 254529 290773 254839 290807
rect 254529 290745 254577 290773
rect 254605 290745 254639 290773
rect 254667 290745 254701 290773
rect 254729 290745 254763 290773
rect 254791 290745 254839 290773
rect 254529 281959 254839 290745
rect 254529 281931 254577 281959
rect 254605 281931 254639 281959
rect 254667 281931 254701 281959
rect 254729 281931 254763 281959
rect 254791 281931 254839 281959
rect 254529 281897 254839 281931
rect 254529 281869 254577 281897
rect 254605 281869 254639 281897
rect 254667 281869 254701 281897
rect 254729 281869 254763 281897
rect 254791 281869 254839 281897
rect 254529 281835 254839 281869
rect 254529 281807 254577 281835
rect 254605 281807 254639 281835
rect 254667 281807 254701 281835
rect 254729 281807 254763 281835
rect 254791 281807 254839 281835
rect 254529 281773 254839 281807
rect 254529 281745 254577 281773
rect 254605 281745 254639 281773
rect 254667 281745 254701 281773
rect 254729 281745 254763 281773
rect 254791 281745 254839 281773
rect 254529 272959 254839 281745
rect 254529 272931 254577 272959
rect 254605 272931 254639 272959
rect 254667 272931 254701 272959
rect 254729 272931 254763 272959
rect 254791 272931 254839 272959
rect 254529 272897 254839 272931
rect 254529 272869 254577 272897
rect 254605 272869 254639 272897
rect 254667 272869 254701 272897
rect 254729 272869 254763 272897
rect 254791 272869 254839 272897
rect 254529 272835 254839 272869
rect 254529 272807 254577 272835
rect 254605 272807 254639 272835
rect 254667 272807 254701 272835
rect 254729 272807 254763 272835
rect 254791 272807 254839 272835
rect 254529 272773 254839 272807
rect 254529 272745 254577 272773
rect 254605 272745 254639 272773
rect 254667 272745 254701 272773
rect 254729 272745 254763 272773
rect 254791 272745 254839 272773
rect 254529 263959 254839 272745
rect 254529 263931 254577 263959
rect 254605 263931 254639 263959
rect 254667 263931 254701 263959
rect 254729 263931 254763 263959
rect 254791 263931 254839 263959
rect 254529 263897 254839 263931
rect 254529 263869 254577 263897
rect 254605 263869 254639 263897
rect 254667 263869 254701 263897
rect 254729 263869 254763 263897
rect 254791 263869 254839 263897
rect 254529 263835 254839 263869
rect 254529 263807 254577 263835
rect 254605 263807 254639 263835
rect 254667 263807 254701 263835
rect 254729 263807 254763 263835
rect 254791 263807 254839 263835
rect 254529 263773 254839 263807
rect 254529 263745 254577 263773
rect 254605 263745 254639 263773
rect 254667 263745 254701 263773
rect 254729 263745 254763 263773
rect 254791 263745 254839 263773
rect 254529 254959 254839 263745
rect 256389 299670 256699 299718
rect 256389 299642 256437 299670
rect 256465 299642 256499 299670
rect 256527 299642 256561 299670
rect 256589 299642 256623 299670
rect 256651 299642 256699 299670
rect 256389 299608 256699 299642
rect 256389 299580 256437 299608
rect 256465 299580 256499 299608
rect 256527 299580 256561 299608
rect 256589 299580 256623 299608
rect 256651 299580 256699 299608
rect 256389 299546 256699 299580
rect 256389 299518 256437 299546
rect 256465 299518 256499 299546
rect 256527 299518 256561 299546
rect 256589 299518 256623 299546
rect 256651 299518 256699 299546
rect 256389 299484 256699 299518
rect 256389 299456 256437 299484
rect 256465 299456 256499 299484
rect 256527 299456 256561 299484
rect 256589 299456 256623 299484
rect 256651 299456 256699 299484
rect 256389 293959 256699 299456
rect 256389 293931 256437 293959
rect 256465 293931 256499 293959
rect 256527 293931 256561 293959
rect 256589 293931 256623 293959
rect 256651 293931 256699 293959
rect 256389 293897 256699 293931
rect 256389 293869 256437 293897
rect 256465 293869 256499 293897
rect 256527 293869 256561 293897
rect 256589 293869 256623 293897
rect 256651 293869 256699 293897
rect 256389 293835 256699 293869
rect 256389 293807 256437 293835
rect 256465 293807 256499 293835
rect 256527 293807 256561 293835
rect 256589 293807 256623 293835
rect 256651 293807 256699 293835
rect 256389 293773 256699 293807
rect 256389 293745 256437 293773
rect 256465 293745 256499 293773
rect 256527 293745 256561 293773
rect 256589 293745 256623 293773
rect 256651 293745 256699 293773
rect 256389 284959 256699 293745
rect 256389 284931 256437 284959
rect 256465 284931 256499 284959
rect 256527 284931 256561 284959
rect 256589 284931 256623 284959
rect 256651 284931 256699 284959
rect 256389 284897 256699 284931
rect 256389 284869 256437 284897
rect 256465 284869 256499 284897
rect 256527 284869 256561 284897
rect 256589 284869 256623 284897
rect 256651 284869 256699 284897
rect 256389 284835 256699 284869
rect 256389 284807 256437 284835
rect 256465 284807 256499 284835
rect 256527 284807 256561 284835
rect 256589 284807 256623 284835
rect 256651 284807 256699 284835
rect 256389 284773 256699 284807
rect 256389 284745 256437 284773
rect 256465 284745 256499 284773
rect 256527 284745 256561 284773
rect 256589 284745 256623 284773
rect 256651 284745 256699 284773
rect 256389 275959 256699 284745
rect 256389 275931 256437 275959
rect 256465 275931 256499 275959
rect 256527 275931 256561 275959
rect 256589 275931 256623 275959
rect 256651 275931 256699 275959
rect 256389 275897 256699 275931
rect 256389 275869 256437 275897
rect 256465 275869 256499 275897
rect 256527 275869 256561 275897
rect 256589 275869 256623 275897
rect 256651 275869 256699 275897
rect 256389 275835 256699 275869
rect 256389 275807 256437 275835
rect 256465 275807 256499 275835
rect 256527 275807 256561 275835
rect 256589 275807 256623 275835
rect 256651 275807 256699 275835
rect 256389 275773 256699 275807
rect 256389 275745 256437 275773
rect 256465 275745 256499 275773
rect 256527 275745 256561 275773
rect 256589 275745 256623 275773
rect 256651 275745 256699 275773
rect 256389 266959 256699 275745
rect 256389 266931 256437 266959
rect 256465 266931 256499 266959
rect 256527 266931 256561 266959
rect 256589 266931 256623 266959
rect 256651 266931 256699 266959
rect 256389 266897 256699 266931
rect 256389 266869 256437 266897
rect 256465 266869 256499 266897
rect 256527 266869 256561 266897
rect 256589 266869 256623 266897
rect 256651 266869 256699 266897
rect 256389 266835 256699 266869
rect 256389 266807 256437 266835
rect 256465 266807 256499 266835
rect 256527 266807 256561 266835
rect 256589 266807 256623 266835
rect 256651 266807 256699 266835
rect 256389 266773 256699 266807
rect 256389 266745 256437 266773
rect 256465 266745 256499 266773
rect 256527 266745 256561 266773
rect 256589 266745 256623 266773
rect 256651 266745 256699 266773
rect 256389 257959 256699 266745
rect 256389 257931 256437 257959
rect 256465 257931 256499 257959
rect 256527 257931 256561 257959
rect 256589 257931 256623 257959
rect 256651 257931 256699 257959
rect 256389 257897 256699 257931
rect 256389 257869 256437 257897
rect 256465 257869 256499 257897
rect 256527 257869 256561 257897
rect 256589 257869 256623 257897
rect 256651 257869 256699 257897
rect 256389 257835 256699 257869
rect 256389 257807 256437 257835
rect 256465 257807 256499 257835
rect 256527 257807 256561 257835
rect 256589 257807 256623 257835
rect 256651 257807 256699 257835
rect 256389 257773 256699 257807
rect 256389 257745 256437 257773
rect 256465 257745 256499 257773
rect 256527 257745 256561 257773
rect 256589 257745 256623 257773
rect 256651 257745 256699 257773
rect 254529 254931 254577 254959
rect 254605 254931 254639 254959
rect 254667 254931 254701 254959
rect 254729 254931 254763 254959
rect 254791 254931 254839 254959
rect 254529 254897 254839 254931
rect 254529 254869 254577 254897
rect 254605 254869 254639 254897
rect 254667 254869 254701 254897
rect 254729 254869 254763 254897
rect 254791 254869 254839 254897
rect 254529 254835 254839 254869
rect 254529 254807 254577 254835
rect 254605 254807 254639 254835
rect 254667 254807 254701 254835
rect 254729 254807 254763 254835
rect 254791 254807 254839 254835
rect 254529 254773 254839 254807
rect 254529 254745 254577 254773
rect 254605 254745 254639 254773
rect 254667 254745 254701 254773
rect 254729 254745 254763 254773
rect 254791 254745 254839 254773
rect 31389 248931 31437 248959
rect 31465 248931 31499 248959
rect 31527 248931 31561 248959
rect 31589 248931 31623 248959
rect 31651 248931 31699 248959
rect 31389 248897 31699 248931
rect 31389 248869 31437 248897
rect 31465 248869 31499 248897
rect 31527 248869 31561 248897
rect 31589 248869 31623 248897
rect 31651 248869 31699 248897
rect 31389 248835 31699 248869
rect 31389 248807 31437 248835
rect 31465 248807 31499 248835
rect 31527 248807 31561 248835
rect 31589 248807 31623 248835
rect 31651 248807 31699 248835
rect 31389 248773 31699 248807
rect 31389 248745 31437 248773
rect 31465 248745 31499 248773
rect 31527 248745 31561 248773
rect 31589 248745 31623 248773
rect 31651 248745 31699 248773
rect 31389 239959 31699 248745
rect 40264 248959 40424 248976
rect 40264 248931 40299 248959
rect 40327 248931 40361 248959
rect 40389 248931 40424 248959
rect 40264 248897 40424 248931
rect 40264 248869 40299 248897
rect 40327 248869 40361 248897
rect 40389 248869 40424 248897
rect 40264 248835 40424 248869
rect 40264 248807 40299 248835
rect 40327 248807 40361 248835
rect 40389 248807 40424 248835
rect 40264 248773 40424 248807
rect 40264 248745 40299 248773
rect 40327 248745 40361 248773
rect 40389 248745 40424 248773
rect 40264 248728 40424 248745
rect 55624 248959 55784 248976
rect 55624 248931 55659 248959
rect 55687 248931 55721 248959
rect 55749 248931 55784 248959
rect 55624 248897 55784 248931
rect 55624 248869 55659 248897
rect 55687 248869 55721 248897
rect 55749 248869 55784 248897
rect 55624 248835 55784 248869
rect 55624 248807 55659 248835
rect 55687 248807 55721 248835
rect 55749 248807 55784 248835
rect 55624 248773 55784 248807
rect 55624 248745 55659 248773
rect 55687 248745 55721 248773
rect 55749 248745 55784 248773
rect 55624 248728 55784 248745
rect 70984 248959 71144 248976
rect 70984 248931 71019 248959
rect 71047 248931 71081 248959
rect 71109 248931 71144 248959
rect 70984 248897 71144 248931
rect 70984 248869 71019 248897
rect 71047 248869 71081 248897
rect 71109 248869 71144 248897
rect 70984 248835 71144 248869
rect 70984 248807 71019 248835
rect 71047 248807 71081 248835
rect 71109 248807 71144 248835
rect 70984 248773 71144 248807
rect 70984 248745 71019 248773
rect 71047 248745 71081 248773
rect 71109 248745 71144 248773
rect 70984 248728 71144 248745
rect 86344 248959 86504 248976
rect 86344 248931 86379 248959
rect 86407 248931 86441 248959
rect 86469 248931 86504 248959
rect 86344 248897 86504 248931
rect 86344 248869 86379 248897
rect 86407 248869 86441 248897
rect 86469 248869 86504 248897
rect 86344 248835 86504 248869
rect 86344 248807 86379 248835
rect 86407 248807 86441 248835
rect 86469 248807 86504 248835
rect 86344 248773 86504 248807
rect 86344 248745 86379 248773
rect 86407 248745 86441 248773
rect 86469 248745 86504 248773
rect 86344 248728 86504 248745
rect 101704 248959 101864 248976
rect 101704 248931 101739 248959
rect 101767 248931 101801 248959
rect 101829 248931 101864 248959
rect 101704 248897 101864 248931
rect 101704 248869 101739 248897
rect 101767 248869 101801 248897
rect 101829 248869 101864 248897
rect 101704 248835 101864 248869
rect 101704 248807 101739 248835
rect 101767 248807 101801 248835
rect 101829 248807 101864 248835
rect 101704 248773 101864 248807
rect 101704 248745 101739 248773
rect 101767 248745 101801 248773
rect 101829 248745 101864 248773
rect 101704 248728 101864 248745
rect 117064 248959 117224 248976
rect 117064 248931 117099 248959
rect 117127 248931 117161 248959
rect 117189 248931 117224 248959
rect 117064 248897 117224 248931
rect 117064 248869 117099 248897
rect 117127 248869 117161 248897
rect 117189 248869 117224 248897
rect 117064 248835 117224 248869
rect 117064 248807 117099 248835
rect 117127 248807 117161 248835
rect 117189 248807 117224 248835
rect 117064 248773 117224 248807
rect 117064 248745 117099 248773
rect 117127 248745 117161 248773
rect 117189 248745 117224 248773
rect 117064 248728 117224 248745
rect 132424 248959 132584 248976
rect 132424 248931 132459 248959
rect 132487 248931 132521 248959
rect 132549 248931 132584 248959
rect 132424 248897 132584 248931
rect 132424 248869 132459 248897
rect 132487 248869 132521 248897
rect 132549 248869 132584 248897
rect 132424 248835 132584 248869
rect 132424 248807 132459 248835
rect 132487 248807 132521 248835
rect 132549 248807 132584 248835
rect 132424 248773 132584 248807
rect 132424 248745 132459 248773
rect 132487 248745 132521 248773
rect 132549 248745 132584 248773
rect 132424 248728 132584 248745
rect 147784 248959 147944 248976
rect 147784 248931 147819 248959
rect 147847 248931 147881 248959
rect 147909 248931 147944 248959
rect 147784 248897 147944 248931
rect 147784 248869 147819 248897
rect 147847 248869 147881 248897
rect 147909 248869 147944 248897
rect 147784 248835 147944 248869
rect 147784 248807 147819 248835
rect 147847 248807 147881 248835
rect 147909 248807 147944 248835
rect 147784 248773 147944 248807
rect 147784 248745 147819 248773
rect 147847 248745 147881 248773
rect 147909 248745 147944 248773
rect 147784 248728 147944 248745
rect 163144 248959 163304 248976
rect 163144 248931 163179 248959
rect 163207 248931 163241 248959
rect 163269 248931 163304 248959
rect 163144 248897 163304 248931
rect 163144 248869 163179 248897
rect 163207 248869 163241 248897
rect 163269 248869 163304 248897
rect 163144 248835 163304 248869
rect 163144 248807 163179 248835
rect 163207 248807 163241 248835
rect 163269 248807 163304 248835
rect 163144 248773 163304 248807
rect 163144 248745 163179 248773
rect 163207 248745 163241 248773
rect 163269 248745 163304 248773
rect 163144 248728 163304 248745
rect 178504 248959 178664 248976
rect 178504 248931 178539 248959
rect 178567 248931 178601 248959
rect 178629 248931 178664 248959
rect 178504 248897 178664 248931
rect 178504 248869 178539 248897
rect 178567 248869 178601 248897
rect 178629 248869 178664 248897
rect 178504 248835 178664 248869
rect 178504 248807 178539 248835
rect 178567 248807 178601 248835
rect 178629 248807 178664 248835
rect 178504 248773 178664 248807
rect 178504 248745 178539 248773
rect 178567 248745 178601 248773
rect 178629 248745 178664 248773
rect 178504 248728 178664 248745
rect 193864 248959 194024 248976
rect 193864 248931 193899 248959
rect 193927 248931 193961 248959
rect 193989 248931 194024 248959
rect 193864 248897 194024 248931
rect 193864 248869 193899 248897
rect 193927 248869 193961 248897
rect 193989 248869 194024 248897
rect 193864 248835 194024 248869
rect 193864 248807 193899 248835
rect 193927 248807 193961 248835
rect 193989 248807 194024 248835
rect 193864 248773 194024 248807
rect 193864 248745 193899 248773
rect 193927 248745 193961 248773
rect 193989 248745 194024 248773
rect 193864 248728 194024 248745
rect 209224 248959 209384 248976
rect 209224 248931 209259 248959
rect 209287 248931 209321 248959
rect 209349 248931 209384 248959
rect 209224 248897 209384 248931
rect 209224 248869 209259 248897
rect 209287 248869 209321 248897
rect 209349 248869 209384 248897
rect 209224 248835 209384 248869
rect 209224 248807 209259 248835
rect 209287 248807 209321 248835
rect 209349 248807 209384 248835
rect 209224 248773 209384 248807
rect 209224 248745 209259 248773
rect 209287 248745 209321 248773
rect 209349 248745 209384 248773
rect 209224 248728 209384 248745
rect 224584 248959 224744 248976
rect 224584 248931 224619 248959
rect 224647 248931 224681 248959
rect 224709 248931 224744 248959
rect 224584 248897 224744 248931
rect 224584 248869 224619 248897
rect 224647 248869 224681 248897
rect 224709 248869 224744 248897
rect 224584 248835 224744 248869
rect 224584 248807 224619 248835
rect 224647 248807 224681 248835
rect 224709 248807 224744 248835
rect 224584 248773 224744 248807
rect 224584 248745 224619 248773
rect 224647 248745 224681 248773
rect 224709 248745 224744 248773
rect 224584 248728 224744 248745
rect 239944 248959 240104 248976
rect 239944 248931 239979 248959
rect 240007 248931 240041 248959
rect 240069 248931 240104 248959
rect 239944 248897 240104 248931
rect 239944 248869 239979 248897
rect 240007 248869 240041 248897
rect 240069 248869 240104 248897
rect 239944 248835 240104 248869
rect 239944 248807 239979 248835
rect 240007 248807 240041 248835
rect 240069 248807 240104 248835
rect 239944 248773 240104 248807
rect 239944 248745 239979 248773
rect 240007 248745 240041 248773
rect 240069 248745 240104 248773
rect 239944 248728 240104 248745
rect 32584 245959 32744 245976
rect 32584 245931 32619 245959
rect 32647 245931 32681 245959
rect 32709 245931 32744 245959
rect 32584 245897 32744 245931
rect 32584 245869 32619 245897
rect 32647 245869 32681 245897
rect 32709 245869 32744 245897
rect 32584 245835 32744 245869
rect 32584 245807 32619 245835
rect 32647 245807 32681 245835
rect 32709 245807 32744 245835
rect 32584 245773 32744 245807
rect 32584 245745 32619 245773
rect 32647 245745 32681 245773
rect 32709 245745 32744 245773
rect 32584 245728 32744 245745
rect 47944 245959 48104 245976
rect 47944 245931 47979 245959
rect 48007 245931 48041 245959
rect 48069 245931 48104 245959
rect 47944 245897 48104 245931
rect 47944 245869 47979 245897
rect 48007 245869 48041 245897
rect 48069 245869 48104 245897
rect 47944 245835 48104 245869
rect 47944 245807 47979 245835
rect 48007 245807 48041 245835
rect 48069 245807 48104 245835
rect 47944 245773 48104 245807
rect 47944 245745 47979 245773
rect 48007 245745 48041 245773
rect 48069 245745 48104 245773
rect 47944 245728 48104 245745
rect 63304 245959 63464 245976
rect 63304 245931 63339 245959
rect 63367 245931 63401 245959
rect 63429 245931 63464 245959
rect 63304 245897 63464 245931
rect 63304 245869 63339 245897
rect 63367 245869 63401 245897
rect 63429 245869 63464 245897
rect 63304 245835 63464 245869
rect 63304 245807 63339 245835
rect 63367 245807 63401 245835
rect 63429 245807 63464 245835
rect 63304 245773 63464 245807
rect 63304 245745 63339 245773
rect 63367 245745 63401 245773
rect 63429 245745 63464 245773
rect 63304 245728 63464 245745
rect 78664 245959 78824 245976
rect 78664 245931 78699 245959
rect 78727 245931 78761 245959
rect 78789 245931 78824 245959
rect 78664 245897 78824 245931
rect 78664 245869 78699 245897
rect 78727 245869 78761 245897
rect 78789 245869 78824 245897
rect 78664 245835 78824 245869
rect 78664 245807 78699 245835
rect 78727 245807 78761 245835
rect 78789 245807 78824 245835
rect 78664 245773 78824 245807
rect 78664 245745 78699 245773
rect 78727 245745 78761 245773
rect 78789 245745 78824 245773
rect 78664 245728 78824 245745
rect 94024 245959 94184 245976
rect 94024 245931 94059 245959
rect 94087 245931 94121 245959
rect 94149 245931 94184 245959
rect 94024 245897 94184 245931
rect 94024 245869 94059 245897
rect 94087 245869 94121 245897
rect 94149 245869 94184 245897
rect 94024 245835 94184 245869
rect 94024 245807 94059 245835
rect 94087 245807 94121 245835
rect 94149 245807 94184 245835
rect 94024 245773 94184 245807
rect 94024 245745 94059 245773
rect 94087 245745 94121 245773
rect 94149 245745 94184 245773
rect 94024 245728 94184 245745
rect 109384 245959 109544 245976
rect 109384 245931 109419 245959
rect 109447 245931 109481 245959
rect 109509 245931 109544 245959
rect 109384 245897 109544 245931
rect 109384 245869 109419 245897
rect 109447 245869 109481 245897
rect 109509 245869 109544 245897
rect 109384 245835 109544 245869
rect 109384 245807 109419 245835
rect 109447 245807 109481 245835
rect 109509 245807 109544 245835
rect 109384 245773 109544 245807
rect 109384 245745 109419 245773
rect 109447 245745 109481 245773
rect 109509 245745 109544 245773
rect 109384 245728 109544 245745
rect 124744 245959 124904 245976
rect 124744 245931 124779 245959
rect 124807 245931 124841 245959
rect 124869 245931 124904 245959
rect 124744 245897 124904 245931
rect 124744 245869 124779 245897
rect 124807 245869 124841 245897
rect 124869 245869 124904 245897
rect 124744 245835 124904 245869
rect 124744 245807 124779 245835
rect 124807 245807 124841 245835
rect 124869 245807 124904 245835
rect 124744 245773 124904 245807
rect 124744 245745 124779 245773
rect 124807 245745 124841 245773
rect 124869 245745 124904 245773
rect 124744 245728 124904 245745
rect 140104 245959 140264 245976
rect 140104 245931 140139 245959
rect 140167 245931 140201 245959
rect 140229 245931 140264 245959
rect 140104 245897 140264 245931
rect 140104 245869 140139 245897
rect 140167 245869 140201 245897
rect 140229 245869 140264 245897
rect 140104 245835 140264 245869
rect 140104 245807 140139 245835
rect 140167 245807 140201 245835
rect 140229 245807 140264 245835
rect 140104 245773 140264 245807
rect 140104 245745 140139 245773
rect 140167 245745 140201 245773
rect 140229 245745 140264 245773
rect 140104 245728 140264 245745
rect 155464 245959 155624 245976
rect 155464 245931 155499 245959
rect 155527 245931 155561 245959
rect 155589 245931 155624 245959
rect 155464 245897 155624 245931
rect 155464 245869 155499 245897
rect 155527 245869 155561 245897
rect 155589 245869 155624 245897
rect 155464 245835 155624 245869
rect 155464 245807 155499 245835
rect 155527 245807 155561 245835
rect 155589 245807 155624 245835
rect 155464 245773 155624 245807
rect 155464 245745 155499 245773
rect 155527 245745 155561 245773
rect 155589 245745 155624 245773
rect 155464 245728 155624 245745
rect 170824 245959 170984 245976
rect 170824 245931 170859 245959
rect 170887 245931 170921 245959
rect 170949 245931 170984 245959
rect 170824 245897 170984 245931
rect 170824 245869 170859 245897
rect 170887 245869 170921 245897
rect 170949 245869 170984 245897
rect 170824 245835 170984 245869
rect 170824 245807 170859 245835
rect 170887 245807 170921 245835
rect 170949 245807 170984 245835
rect 170824 245773 170984 245807
rect 170824 245745 170859 245773
rect 170887 245745 170921 245773
rect 170949 245745 170984 245773
rect 170824 245728 170984 245745
rect 186184 245959 186344 245976
rect 186184 245931 186219 245959
rect 186247 245931 186281 245959
rect 186309 245931 186344 245959
rect 186184 245897 186344 245931
rect 186184 245869 186219 245897
rect 186247 245869 186281 245897
rect 186309 245869 186344 245897
rect 186184 245835 186344 245869
rect 186184 245807 186219 245835
rect 186247 245807 186281 245835
rect 186309 245807 186344 245835
rect 186184 245773 186344 245807
rect 186184 245745 186219 245773
rect 186247 245745 186281 245773
rect 186309 245745 186344 245773
rect 186184 245728 186344 245745
rect 201544 245959 201704 245976
rect 201544 245931 201579 245959
rect 201607 245931 201641 245959
rect 201669 245931 201704 245959
rect 201544 245897 201704 245931
rect 201544 245869 201579 245897
rect 201607 245869 201641 245897
rect 201669 245869 201704 245897
rect 201544 245835 201704 245869
rect 201544 245807 201579 245835
rect 201607 245807 201641 245835
rect 201669 245807 201704 245835
rect 201544 245773 201704 245807
rect 201544 245745 201579 245773
rect 201607 245745 201641 245773
rect 201669 245745 201704 245773
rect 201544 245728 201704 245745
rect 216904 245959 217064 245976
rect 216904 245931 216939 245959
rect 216967 245931 217001 245959
rect 217029 245931 217064 245959
rect 216904 245897 217064 245931
rect 216904 245869 216939 245897
rect 216967 245869 217001 245897
rect 217029 245869 217064 245897
rect 216904 245835 217064 245869
rect 216904 245807 216939 245835
rect 216967 245807 217001 245835
rect 217029 245807 217064 245835
rect 216904 245773 217064 245807
rect 216904 245745 216939 245773
rect 216967 245745 217001 245773
rect 217029 245745 217064 245773
rect 216904 245728 217064 245745
rect 232264 245959 232424 245976
rect 232264 245931 232299 245959
rect 232327 245931 232361 245959
rect 232389 245931 232424 245959
rect 232264 245897 232424 245931
rect 232264 245869 232299 245897
rect 232327 245869 232361 245897
rect 232389 245869 232424 245897
rect 232264 245835 232424 245869
rect 232264 245807 232299 245835
rect 232327 245807 232361 245835
rect 232389 245807 232424 245835
rect 232264 245773 232424 245807
rect 232264 245745 232299 245773
rect 232327 245745 232361 245773
rect 232389 245745 232424 245773
rect 232264 245728 232424 245745
rect 247624 245959 247784 245976
rect 247624 245931 247659 245959
rect 247687 245931 247721 245959
rect 247749 245931 247784 245959
rect 247624 245897 247784 245931
rect 247624 245869 247659 245897
rect 247687 245869 247721 245897
rect 247749 245869 247784 245897
rect 247624 245835 247784 245869
rect 247624 245807 247659 245835
rect 247687 245807 247721 245835
rect 247749 245807 247784 245835
rect 247624 245773 247784 245807
rect 247624 245745 247659 245773
rect 247687 245745 247721 245773
rect 247749 245745 247784 245773
rect 247624 245728 247784 245745
rect 254529 245959 254839 254745
rect 254529 245931 254577 245959
rect 254605 245931 254639 245959
rect 254667 245931 254701 245959
rect 254729 245931 254763 245959
rect 254791 245931 254839 245959
rect 254529 245897 254839 245931
rect 254529 245869 254577 245897
rect 254605 245869 254639 245897
rect 254667 245869 254701 245897
rect 254729 245869 254763 245897
rect 254791 245869 254839 245897
rect 254529 245835 254839 245869
rect 254529 245807 254577 245835
rect 254605 245807 254639 245835
rect 254667 245807 254701 245835
rect 254729 245807 254763 245835
rect 254791 245807 254839 245835
rect 254529 245773 254839 245807
rect 254529 245745 254577 245773
rect 254605 245745 254639 245773
rect 254667 245745 254701 245773
rect 254729 245745 254763 245773
rect 254791 245745 254839 245773
rect 31389 239931 31437 239959
rect 31465 239931 31499 239959
rect 31527 239931 31561 239959
rect 31589 239931 31623 239959
rect 31651 239931 31699 239959
rect 31389 239897 31699 239931
rect 31389 239869 31437 239897
rect 31465 239869 31499 239897
rect 31527 239869 31561 239897
rect 31589 239869 31623 239897
rect 31651 239869 31699 239897
rect 31389 239835 31699 239869
rect 31389 239807 31437 239835
rect 31465 239807 31499 239835
rect 31527 239807 31561 239835
rect 31589 239807 31623 239835
rect 31651 239807 31699 239835
rect 31389 239773 31699 239807
rect 31389 239745 31437 239773
rect 31465 239745 31499 239773
rect 31527 239745 31561 239773
rect 31589 239745 31623 239773
rect 31651 239745 31699 239773
rect 31389 230959 31699 239745
rect 40264 239959 40424 239976
rect 40264 239931 40299 239959
rect 40327 239931 40361 239959
rect 40389 239931 40424 239959
rect 40264 239897 40424 239931
rect 40264 239869 40299 239897
rect 40327 239869 40361 239897
rect 40389 239869 40424 239897
rect 40264 239835 40424 239869
rect 40264 239807 40299 239835
rect 40327 239807 40361 239835
rect 40389 239807 40424 239835
rect 40264 239773 40424 239807
rect 40264 239745 40299 239773
rect 40327 239745 40361 239773
rect 40389 239745 40424 239773
rect 40264 239728 40424 239745
rect 55624 239959 55784 239976
rect 55624 239931 55659 239959
rect 55687 239931 55721 239959
rect 55749 239931 55784 239959
rect 55624 239897 55784 239931
rect 55624 239869 55659 239897
rect 55687 239869 55721 239897
rect 55749 239869 55784 239897
rect 55624 239835 55784 239869
rect 55624 239807 55659 239835
rect 55687 239807 55721 239835
rect 55749 239807 55784 239835
rect 55624 239773 55784 239807
rect 55624 239745 55659 239773
rect 55687 239745 55721 239773
rect 55749 239745 55784 239773
rect 55624 239728 55784 239745
rect 70984 239959 71144 239976
rect 70984 239931 71019 239959
rect 71047 239931 71081 239959
rect 71109 239931 71144 239959
rect 70984 239897 71144 239931
rect 70984 239869 71019 239897
rect 71047 239869 71081 239897
rect 71109 239869 71144 239897
rect 70984 239835 71144 239869
rect 70984 239807 71019 239835
rect 71047 239807 71081 239835
rect 71109 239807 71144 239835
rect 70984 239773 71144 239807
rect 70984 239745 71019 239773
rect 71047 239745 71081 239773
rect 71109 239745 71144 239773
rect 70984 239728 71144 239745
rect 86344 239959 86504 239976
rect 86344 239931 86379 239959
rect 86407 239931 86441 239959
rect 86469 239931 86504 239959
rect 86344 239897 86504 239931
rect 86344 239869 86379 239897
rect 86407 239869 86441 239897
rect 86469 239869 86504 239897
rect 86344 239835 86504 239869
rect 86344 239807 86379 239835
rect 86407 239807 86441 239835
rect 86469 239807 86504 239835
rect 86344 239773 86504 239807
rect 86344 239745 86379 239773
rect 86407 239745 86441 239773
rect 86469 239745 86504 239773
rect 86344 239728 86504 239745
rect 101704 239959 101864 239976
rect 101704 239931 101739 239959
rect 101767 239931 101801 239959
rect 101829 239931 101864 239959
rect 101704 239897 101864 239931
rect 101704 239869 101739 239897
rect 101767 239869 101801 239897
rect 101829 239869 101864 239897
rect 101704 239835 101864 239869
rect 101704 239807 101739 239835
rect 101767 239807 101801 239835
rect 101829 239807 101864 239835
rect 101704 239773 101864 239807
rect 101704 239745 101739 239773
rect 101767 239745 101801 239773
rect 101829 239745 101864 239773
rect 101704 239728 101864 239745
rect 117064 239959 117224 239976
rect 117064 239931 117099 239959
rect 117127 239931 117161 239959
rect 117189 239931 117224 239959
rect 117064 239897 117224 239931
rect 117064 239869 117099 239897
rect 117127 239869 117161 239897
rect 117189 239869 117224 239897
rect 117064 239835 117224 239869
rect 117064 239807 117099 239835
rect 117127 239807 117161 239835
rect 117189 239807 117224 239835
rect 117064 239773 117224 239807
rect 117064 239745 117099 239773
rect 117127 239745 117161 239773
rect 117189 239745 117224 239773
rect 117064 239728 117224 239745
rect 132424 239959 132584 239976
rect 132424 239931 132459 239959
rect 132487 239931 132521 239959
rect 132549 239931 132584 239959
rect 132424 239897 132584 239931
rect 132424 239869 132459 239897
rect 132487 239869 132521 239897
rect 132549 239869 132584 239897
rect 132424 239835 132584 239869
rect 132424 239807 132459 239835
rect 132487 239807 132521 239835
rect 132549 239807 132584 239835
rect 132424 239773 132584 239807
rect 132424 239745 132459 239773
rect 132487 239745 132521 239773
rect 132549 239745 132584 239773
rect 132424 239728 132584 239745
rect 147784 239959 147944 239976
rect 147784 239931 147819 239959
rect 147847 239931 147881 239959
rect 147909 239931 147944 239959
rect 147784 239897 147944 239931
rect 147784 239869 147819 239897
rect 147847 239869 147881 239897
rect 147909 239869 147944 239897
rect 147784 239835 147944 239869
rect 147784 239807 147819 239835
rect 147847 239807 147881 239835
rect 147909 239807 147944 239835
rect 147784 239773 147944 239807
rect 147784 239745 147819 239773
rect 147847 239745 147881 239773
rect 147909 239745 147944 239773
rect 147784 239728 147944 239745
rect 163144 239959 163304 239976
rect 163144 239931 163179 239959
rect 163207 239931 163241 239959
rect 163269 239931 163304 239959
rect 163144 239897 163304 239931
rect 163144 239869 163179 239897
rect 163207 239869 163241 239897
rect 163269 239869 163304 239897
rect 163144 239835 163304 239869
rect 163144 239807 163179 239835
rect 163207 239807 163241 239835
rect 163269 239807 163304 239835
rect 163144 239773 163304 239807
rect 163144 239745 163179 239773
rect 163207 239745 163241 239773
rect 163269 239745 163304 239773
rect 163144 239728 163304 239745
rect 178504 239959 178664 239976
rect 178504 239931 178539 239959
rect 178567 239931 178601 239959
rect 178629 239931 178664 239959
rect 178504 239897 178664 239931
rect 178504 239869 178539 239897
rect 178567 239869 178601 239897
rect 178629 239869 178664 239897
rect 178504 239835 178664 239869
rect 178504 239807 178539 239835
rect 178567 239807 178601 239835
rect 178629 239807 178664 239835
rect 178504 239773 178664 239807
rect 178504 239745 178539 239773
rect 178567 239745 178601 239773
rect 178629 239745 178664 239773
rect 178504 239728 178664 239745
rect 193864 239959 194024 239976
rect 193864 239931 193899 239959
rect 193927 239931 193961 239959
rect 193989 239931 194024 239959
rect 193864 239897 194024 239931
rect 193864 239869 193899 239897
rect 193927 239869 193961 239897
rect 193989 239869 194024 239897
rect 193864 239835 194024 239869
rect 193864 239807 193899 239835
rect 193927 239807 193961 239835
rect 193989 239807 194024 239835
rect 193864 239773 194024 239807
rect 193864 239745 193899 239773
rect 193927 239745 193961 239773
rect 193989 239745 194024 239773
rect 193864 239728 194024 239745
rect 209224 239959 209384 239976
rect 209224 239931 209259 239959
rect 209287 239931 209321 239959
rect 209349 239931 209384 239959
rect 209224 239897 209384 239931
rect 209224 239869 209259 239897
rect 209287 239869 209321 239897
rect 209349 239869 209384 239897
rect 209224 239835 209384 239869
rect 209224 239807 209259 239835
rect 209287 239807 209321 239835
rect 209349 239807 209384 239835
rect 209224 239773 209384 239807
rect 209224 239745 209259 239773
rect 209287 239745 209321 239773
rect 209349 239745 209384 239773
rect 209224 239728 209384 239745
rect 224584 239959 224744 239976
rect 224584 239931 224619 239959
rect 224647 239931 224681 239959
rect 224709 239931 224744 239959
rect 224584 239897 224744 239931
rect 224584 239869 224619 239897
rect 224647 239869 224681 239897
rect 224709 239869 224744 239897
rect 224584 239835 224744 239869
rect 224584 239807 224619 239835
rect 224647 239807 224681 239835
rect 224709 239807 224744 239835
rect 224584 239773 224744 239807
rect 224584 239745 224619 239773
rect 224647 239745 224681 239773
rect 224709 239745 224744 239773
rect 224584 239728 224744 239745
rect 239944 239959 240104 239976
rect 239944 239931 239979 239959
rect 240007 239931 240041 239959
rect 240069 239931 240104 239959
rect 239944 239897 240104 239931
rect 239944 239869 239979 239897
rect 240007 239869 240041 239897
rect 240069 239869 240104 239897
rect 239944 239835 240104 239869
rect 239944 239807 239979 239835
rect 240007 239807 240041 239835
rect 240069 239807 240104 239835
rect 239944 239773 240104 239807
rect 239944 239745 239979 239773
rect 240007 239745 240041 239773
rect 240069 239745 240104 239773
rect 239944 239728 240104 239745
rect 32584 236959 32744 236976
rect 32584 236931 32619 236959
rect 32647 236931 32681 236959
rect 32709 236931 32744 236959
rect 32584 236897 32744 236931
rect 32584 236869 32619 236897
rect 32647 236869 32681 236897
rect 32709 236869 32744 236897
rect 32584 236835 32744 236869
rect 32584 236807 32619 236835
rect 32647 236807 32681 236835
rect 32709 236807 32744 236835
rect 32584 236773 32744 236807
rect 32584 236745 32619 236773
rect 32647 236745 32681 236773
rect 32709 236745 32744 236773
rect 32584 236728 32744 236745
rect 47944 236959 48104 236976
rect 47944 236931 47979 236959
rect 48007 236931 48041 236959
rect 48069 236931 48104 236959
rect 47944 236897 48104 236931
rect 47944 236869 47979 236897
rect 48007 236869 48041 236897
rect 48069 236869 48104 236897
rect 47944 236835 48104 236869
rect 47944 236807 47979 236835
rect 48007 236807 48041 236835
rect 48069 236807 48104 236835
rect 47944 236773 48104 236807
rect 47944 236745 47979 236773
rect 48007 236745 48041 236773
rect 48069 236745 48104 236773
rect 47944 236728 48104 236745
rect 63304 236959 63464 236976
rect 63304 236931 63339 236959
rect 63367 236931 63401 236959
rect 63429 236931 63464 236959
rect 63304 236897 63464 236931
rect 63304 236869 63339 236897
rect 63367 236869 63401 236897
rect 63429 236869 63464 236897
rect 63304 236835 63464 236869
rect 63304 236807 63339 236835
rect 63367 236807 63401 236835
rect 63429 236807 63464 236835
rect 63304 236773 63464 236807
rect 63304 236745 63339 236773
rect 63367 236745 63401 236773
rect 63429 236745 63464 236773
rect 63304 236728 63464 236745
rect 78664 236959 78824 236976
rect 78664 236931 78699 236959
rect 78727 236931 78761 236959
rect 78789 236931 78824 236959
rect 78664 236897 78824 236931
rect 78664 236869 78699 236897
rect 78727 236869 78761 236897
rect 78789 236869 78824 236897
rect 78664 236835 78824 236869
rect 78664 236807 78699 236835
rect 78727 236807 78761 236835
rect 78789 236807 78824 236835
rect 78664 236773 78824 236807
rect 78664 236745 78699 236773
rect 78727 236745 78761 236773
rect 78789 236745 78824 236773
rect 78664 236728 78824 236745
rect 94024 236959 94184 236976
rect 94024 236931 94059 236959
rect 94087 236931 94121 236959
rect 94149 236931 94184 236959
rect 94024 236897 94184 236931
rect 94024 236869 94059 236897
rect 94087 236869 94121 236897
rect 94149 236869 94184 236897
rect 94024 236835 94184 236869
rect 94024 236807 94059 236835
rect 94087 236807 94121 236835
rect 94149 236807 94184 236835
rect 94024 236773 94184 236807
rect 94024 236745 94059 236773
rect 94087 236745 94121 236773
rect 94149 236745 94184 236773
rect 94024 236728 94184 236745
rect 109384 236959 109544 236976
rect 109384 236931 109419 236959
rect 109447 236931 109481 236959
rect 109509 236931 109544 236959
rect 109384 236897 109544 236931
rect 109384 236869 109419 236897
rect 109447 236869 109481 236897
rect 109509 236869 109544 236897
rect 109384 236835 109544 236869
rect 109384 236807 109419 236835
rect 109447 236807 109481 236835
rect 109509 236807 109544 236835
rect 109384 236773 109544 236807
rect 109384 236745 109419 236773
rect 109447 236745 109481 236773
rect 109509 236745 109544 236773
rect 109384 236728 109544 236745
rect 124744 236959 124904 236976
rect 124744 236931 124779 236959
rect 124807 236931 124841 236959
rect 124869 236931 124904 236959
rect 124744 236897 124904 236931
rect 124744 236869 124779 236897
rect 124807 236869 124841 236897
rect 124869 236869 124904 236897
rect 124744 236835 124904 236869
rect 124744 236807 124779 236835
rect 124807 236807 124841 236835
rect 124869 236807 124904 236835
rect 124744 236773 124904 236807
rect 124744 236745 124779 236773
rect 124807 236745 124841 236773
rect 124869 236745 124904 236773
rect 124744 236728 124904 236745
rect 140104 236959 140264 236976
rect 140104 236931 140139 236959
rect 140167 236931 140201 236959
rect 140229 236931 140264 236959
rect 140104 236897 140264 236931
rect 140104 236869 140139 236897
rect 140167 236869 140201 236897
rect 140229 236869 140264 236897
rect 140104 236835 140264 236869
rect 140104 236807 140139 236835
rect 140167 236807 140201 236835
rect 140229 236807 140264 236835
rect 140104 236773 140264 236807
rect 140104 236745 140139 236773
rect 140167 236745 140201 236773
rect 140229 236745 140264 236773
rect 140104 236728 140264 236745
rect 155464 236959 155624 236976
rect 155464 236931 155499 236959
rect 155527 236931 155561 236959
rect 155589 236931 155624 236959
rect 155464 236897 155624 236931
rect 155464 236869 155499 236897
rect 155527 236869 155561 236897
rect 155589 236869 155624 236897
rect 155464 236835 155624 236869
rect 155464 236807 155499 236835
rect 155527 236807 155561 236835
rect 155589 236807 155624 236835
rect 155464 236773 155624 236807
rect 155464 236745 155499 236773
rect 155527 236745 155561 236773
rect 155589 236745 155624 236773
rect 155464 236728 155624 236745
rect 170824 236959 170984 236976
rect 170824 236931 170859 236959
rect 170887 236931 170921 236959
rect 170949 236931 170984 236959
rect 170824 236897 170984 236931
rect 170824 236869 170859 236897
rect 170887 236869 170921 236897
rect 170949 236869 170984 236897
rect 170824 236835 170984 236869
rect 170824 236807 170859 236835
rect 170887 236807 170921 236835
rect 170949 236807 170984 236835
rect 170824 236773 170984 236807
rect 170824 236745 170859 236773
rect 170887 236745 170921 236773
rect 170949 236745 170984 236773
rect 170824 236728 170984 236745
rect 186184 236959 186344 236976
rect 186184 236931 186219 236959
rect 186247 236931 186281 236959
rect 186309 236931 186344 236959
rect 186184 236897 186344 236931
rect 186184 236869 186219 236897
rect 186247 236869 186281 236897
rect 186309 236869 186344 236897
rect 186184 236835 186344 236869
rect 186184 236807 186219 236835
rect 186247 236807 186281 236835
rect 186309 236807 186344 236835
rect 186184 236773 186344 236807
rect 186184 236745 186219 236773
rect 186247 236745 186281 236773
rect 186309 236745 186344 236773
rect 186184 236728 186344 236745
rect 201544 236959 201704 236976
rect 201544 236931 201579 236959
rect 201607 236931 201641 236959
rect 201669 236931 201704 236959
rect 201544 236897 201704 236931
rect 201544 236869 201579 236897
rect 201607 236869 201641 236897
rect 201669 236869 201704 236897
rect 201544 236835 201704 236869
rect 201544 236807 201579 236835
rect 201607 236807 201641 236835
rect 201669 236807 201704 236835
rect 201544 236773 201704 236807
rect 201544 236745 201579 236773
rect 201607 236745 201641 236773
rect 201669 236745 201704 236773
rect 201544 236728 201704 236745
rect 216904 236959 217064 236976
rect 216904 236931 216939 236959
rect 216967 236931 217001 236959
rect 217029 236931 217064 236959
rect 216904 236897 217064 236931
rect 216904 236869 216939 236897
rect 216967 236869 217001 236897
rect 217029 236869 217064 236897
rect 216904 236835 217064 236869
rect 216904 236807 216939 236835
rect 216967 236807 217001 236835
rect 217029 236807 217064 236835
rect 216904 236773 217064 236807
rect 216904 236745 216939 236773
rect 216967 236745 217001 236773
rect 217029 236745 217064 236773
rect 216904 236728 217064 236745
rect 232264 236959 232424 236976
rect 232264 236931 232299 236959
rect 232327 236931 232361 236959
rect 232389 236931 232424 236959
rect 232264 236897 232424 236931
rect 232264 236869 232299 236897
rect 232327 236869 232361 236897
rect 232389 236869 232424 236897
rect 232264 236835 232424 236869
rect 232264 236807 232299 236835
rect 232327 236807 232361 236835
rect 232389 236807 232424 236835
rect 232264 236773 232424 236807
rect 232264 236745 232299 236773
rect 232327 236745 232361 236773
rect 232389 236745 232424 236773
rect 232264 236728 232424 236745
rect 247624 236959 247784 236976
rect 247624 236931 247659 236959
rect 247687 236931 247721 236959
rect 247749 236931 247784 236959
rect 247624 236897 247784 236931
rect 247624 236869 247659 236897
rect 247687 236869 247721 236897
rect 247749 236869 247784 236897
rect 247624 236835 247784 236869
rect 247624 236807 247659 236835
rect 247687 236807 247721 236835
rect 247749 236807 247784 236835
rect 247624 236773 247784 236807
rect 247624 236745 247659 236773
rect 247687 236745 247721 236773
rect 247749 236745 247784 236773
rect 247624 236728 247784 236745
rect 254529 236959 254839 245745
rect 254529 236931 254577 236959
rect 254605 236931 254639 236959
rect 254667 236931 254701 236959
rect 254729 236931 254763 236959
rect 254791 236931 254839 236959
rect 254529 236897 254839 236931
rect 254529 236869 254577 236897
rect 254605 236869 254639 236897
rect 254667 236869 254701 236897
rect 254729 236869 254763 236897
rect 254791 236869 254839 236897
rect 254529 236835 254839 236869
rect 254529 236807 254577 236835
rect 254605 236807 254639 236835
rect 254667 236807 254701 236835
rect 254729 236807 254763 236835
rect 254791 236807 254839 236835
rect 254529 236773 254839 236807
rect 254529 236745 254577 236773
rect 254605 236745 254639 236773
rect 254667 236745 254701 236773
rect 254729 236745 254763 236773
rect 254791 236745 254839 236773
rect 31389 230931 31437 230959
rect 31465 230931 31499 230959
rect 31527 230931 31561 230959
rect 31589 230931 31623 230959
rect 31651 230931 31699 230959
rect 31389 230897 31699 230931
rect 31389 230869 31437 230897
rect 31465 230869 31499 230897
rect 31527 230869 31561 230897
rect 31589 230869 31623 230897
rect 31651 230869 31699 230897
rect 31389 230835 31699 230869
rect 31389 230807 31437 230835
rect 31465 230807 31499 230835
rect 31527 230807 31561 230835
rect 31589 230807 31623 230835
rect 31651 230807 31699 230835
rect 31389 230773 31699 230807
rect 31389 230745 31437 230773
rect 31465 230745 31499 230773
rect 31527 230745 31561 230773
rect 31589 230745 31623 230773
rect 31651 230745 31699 230773
rect 31389 221959 31699 230745
rect 40264 230959 40424 230976
rect 40264 230931 40299 230959
rect 40327 230931 40361 230959
rect 40389 230931 40424 230959
rect 40264 230897 40424 230931
rect 40264 230869 40299 230897
rect 40327 230869 40361 230897
rect 40389 230869 40424 230897
rect 40264 230835 40424 230869
rect 40264 230807 40299 230835
rect 40327 230807 40361 230835
rect 40389 230807 40424 230835
rect 40264 230773 40424 230807
rect 40264 230745 40299 230773
rect 40327 230745 40361 230773
rect 40389 230745 40424 230773
rect 40264 230728 40424 230745
rect 55624 230959 55784 230976
rect 55624 230931 55659 230959
rect 55687 230931 55721 230959
rect 55749 230931 55784 230959
rect 55624 230897 55784 230931
rect 55624 230869 55659 230897
rect 55687 230869 55721 230897
rect 55749 230869 55784 230897
rect 55624 230835 55784 230869
rect 55624 230807 55659 230835
rect 55687 230807 55721 230835
rect 55749 230807 55784 230835
rect 55624 230773 55784 230807
rect 55624 230745 55659 230773
rect 55687 230745 55721 230773
rect 55749 230745 55784 230773
rect 55624 230728 55784 230745
rect 70984 230959 71144 230976
rect 70984 230931 71019 230959
rect 71047 230931 71081 230959
rect 71109 230931 71144 230959
rect 70984 230897 71144 230931
rect 70984 230869 71019 230897
rect 71047 230869 71081 230897
rect 71109 230869 71144 230897
rect 70984 230835 71144 230869
rect 70984 230807 71019 230835
rect 71047 230807 71081 230835
rect 71109 230807 71144 230835
rect 70984 230773 71144 230807
rect 70984 230745 71019 230773
rect 71047 230745 71081 230773
rect 71109 230745 71144 230773
rect 70984 230728 71144 230745
rect 86344 230959 86504 230976
rect 86344 230931 86379 230959
rect 86407 230931 86441 230959
rect 86469 230931 86504 230959
rect 86344 230897 86504 230931
rect 86344 230869 86379 230897
rect 86407 230869 86441 230897
rect 86469 230869 86504 230897
rect 86344 230835 86504 230869
rect 86344 230807 86379 230835
rect 86407 230807 86441 230835
rect 86469 230807 86504 230835
rect 86344 230773 86504 230807
rect 86344 230745 86379 230773
rect 86407 230745 86441 230773
rect 86469 230745 86504 230773
rect 86344 230728 86504 230745
rect 101704 230959 101864 230976
rect 101704 230931 101739 230959
rect 101767 230931 101801 230959
rect 101829 230931 101864 230959
rect 101704 230897 101864 230931
rect 101704 230869 101739 230897
rect 101767 230869 101801 230897
rect 101829 230869 101864 230897
rect 101704 230835 101864 230869
rect 101704 230807 101739 230835
rect 101767 230807 101801 230835
rect 101829 230807 101864 230835
rect 101704 230773 101864 230807
rect 101704 230745 101739 230773
rect 101767 230745 101801 230773
rect 101829 230745 101864 230773
rect 101704 230728 101864 230745
rect 117064 230959 117224 230976
rect 117064 230931 117099 230959
rect 117127 230931 117161 230959
rect 117189 230931 117224 230959
rect 117064 230897 117224 230931
rect 117064 230869 117099 230897
rect 117127 230869 117161 230897
rect 117189 230869 117224 230897
rect 117064 230835 117224 230869
rect 117064 230807 117099 230835
rect 117127 230807 117161 230835
rect 117189 230807 117224 230835
rect 117064 230773 117224 230807
rect 117064 230745 117099 230773
rect 117127 230745 117161 230773
rect 117189 230745 117224 230773
rect 117064 230728 117224 230745
rect 132424 230959 132584 230976
rect 132424 230931 132459 230959
rect 132487 230931 132521 230959
rect 132549 230931 132584 230959
rect 132424 230897 132584 230931
rect 132424 230869 132459 230897
rect 132487 230869 132521 230897
rect 132549 230869 132584 230897
rect 132424 230835 132584 230869
rect 132424 230807 132459 230835
rect 132487 230807 132521 230835
rect 132549 230807 132584 230835
rect 132424 230773 132584 230807
rect 132424 230745 132459 230773
rect 132487 230745 132521 230773
rect 132549 230745 132584 230773
rect 132424 230728 132584 230745
rect 147784 230959 147944 230976
rect 147784 230931 147819 230959
rect 147847 230931 147881 230959
rect 147909 230931 147944 230959
rect 147784 230897 147944 230931
rect 147784 230869 147819 230897
rect 147847 230869 147881 230897
rect 147909 230869 147944 230897
rect 147784 230835 147944 230869
rect 147784 230807 147819 230835
rect 147847 230807 147881 230835
rect 147909 230807 147944 230835
rect 147784 230773 147944 230807
rect 147784 230745 147819 230773
rect 147847 230745 147881 230773
rect 147909 230745 147944 230773
rect 147784 230728 147944 230745
rect 163144 230959 163304 230976
rect 163144 230931 163179 230959
rect 163207 230931 163241 230959
rect 163269 230931 163304 230959
rect 163144 230897 163304 230931
rect 163144 230869 163179 230897
rect 163207 230869 163241 230897
rect 163269 230869 163304 230897
rect 163144 230835 163304 230869
rect 163144 230807 163179 230835
rect 163207 230807 163241 230835
rect 163269 230807 163304 230835
rect 163144 230773 163304 230807
rect 163144 230745 163179 230773
rect 163207 230745 163241 230773
rect 163269 230745 163304 230773
rect 163144 230728 163304 230745
rect 178504 230959 178664 230976
rect 178504 230931 178539 230959
rect 178567 230931 178601 230959
rect 178629 230931 178664 230959
rect 178504 230897 178664 230931
rect 178504 230869 178539 230897
rect 178567 230869 178601 230897
rect 178629 230869 178664 230897
rect 178504 230835 178664 230869
rect 178504 230807 178539 230835
rect 178567 230807 178601 230835
rect 178629 230807 178664 230835
rect 178504 230773 178664 230807
rect 178504 230745 178539 230773
rect 178567 230745 178601 230773
rect 178629 230745 178664 230773
rect 178504 230728 178664 230745
rect 193864 230959 194024 230976
rect 193864 230931 193899 230959
rect 193927 230931 193961 230959
rect 193989 230931 194024 230959
rect 193864 230897 194024 230931
rect 193864 230869 193899 230897
rect 193927 230869 193961 230897
rect 193989 230869 194024 230897
rect 193864 230835 194024 230869
rect 193864 230807 193899 230835
rect 193927 230807 193961 230835
rect 193989 230807 194024 230835
rect 193864 230773 194024 230807
rect 193864 230745 193899 230773
rect 193927 230745 193961 230773
rect 193989 230745 194024 230773
rect 193864 230728 194024 230745
rect 209224 230959 209384 230976
rect 209224 230931 209259 230959
rect 209287 230931 209321 230959
rect 209349 230931 209384 230959
rect 209224 230897 209384 230931
rect 209224 230869 209259 230897
rect 209287 230869 209321 230897
rect 209349 230869 209384 230897
rect 209224 230835 209384 230869
rect 209224 230807 209259 230835
rect 209287 230807 209321 230835
rect 209349 230807 209384 230835
rect 209224 230773 209384 230807
rect 209224 230745 209259 230773
rect 209287 230745 209321 230773
rect 209349 230745 209384 230773
rect 209224 230728 209384 230745
rect 224584 230959 224744 230976
rect 224584 230931 224619 230959
rect 224647 230931 224681 230959
rect 224709 230931 224744 230959
rect 224584 230897 224744 230931
rect 224584 230869 224619 230897
rect 224647 230869 224681 230897
rect 224709 230869 224744 230897
rect 224584 230835 224744 230869
rect 224584 230807 224619 230835
rect 224647 230807 224681 230835
rect 224709 230807 224744 230835
rect 224584 230773 224744 230807
rect 224584 230745 224619 230773
rect 224647 230745 224681 230773
rect 224709 230745 224744 230773
rect 224584 230728 224744 230745
rect 239944 230959 240104 230976
rect 239944 230931 239979 230959
rect 240007 230931 240041 230959
rect 240069 230931 240104 230959
rect 239944 230897 240104 230931
rect 239944 230869 239979 230897
rect 240007 230869 240041 230897
rect 240069 230869 240104 230897
rect 239944 230835 240104 230869
rect 239944 230807 239979 230835
rect 240007 230807 240041 230835
rect 240069 230807 240104 230835
rect 239944 230773 240104 230807
rect 239944 230745 239979 230773
rect 240007 230745 240041 230773
rect 240069 230745 240104 230773
rect 239944 230728 240104 230745
rect 32584 227959 32744 227976
rect 32584 227931 32619 227959
rect 32647 227931 32681 227959
rect 32709 227931 32744 227959
rect 32584 227897 32744 227931
rect 32584 227869 32619 227897
rect 32647 227869 32681 227897
rect 32709 227869 32744 227897
rect 32584 227835 32744 227869
rect 32584 227807 32619 227835
rect 32647 227807 32681 227835
rect 32709 227807 32744 227835
rect 32584 227773 32744 227807
rect 32584 227745 32619 227773
rect 32647 227745 32681 227773
rect 32709 227745 32744 227773
rect 32584 227728 32744 227745
rect 47944 227959 48104 227976
rect 47944 227931 47979 227959
rect 48007 227931 48041 227959
rect 48069 227931 48104 227959
rect 47944 227897 48104 227931
rect 47944 227869 47979 227897
rect 48007 227869 48041 227897
rect 48069 227869 48104 227897
rect 47944 227835 48104 227869
rect 47944 227807 47979 227835
rect 48007 227807 48041 227835
rect 48069 227807 48104 227835
rect 47944 227773 48104 227807
rect 47944 227745 47979 227773
rect 48007 227745 48041 227773
rect 48069 227745 48104 227773
rect 47944 227728 48104 227745
rect 63304 227959 63464 227976
rect 63304 227931 63339 227959
rect 63367 227931 63401 227959
rect 63429 227931 63464 227959
rect 63304 227897 63464 227931
rect 63304 227869 63339 227897
rect 63367 227869 63401 227897
rect 63429 227869 63464 227897
rect 63304 227835 63464 227869
rect 63304 227807 63339 227835
rect 63367 227807 63401 227835
rect 63429 227807 63464 227835
rect 63304 227773 63464 227807
rect 63304 227745 63339 227773
rect 63367 227745 63401 227773
rect 63429 227745 63464 227773
rect 63304 227728 63464 227745
rect 78664 227959 78824 227976
rect 78664 227931 78699 227959
rect 78727 227931 78761 227959
rect 78789 227931 78824 227959
rect 78664 227897 78824 227931
rect 78664 227869 78699 227897
rect 78727 227869 78761 227897
rect 78789 227869 78824 227897
rect 78664 227835 78824 227869
rect 78664 227807 78699 227835
rect 78727 227807 78761 227835
rect 78789 227807 78824 227835
rect 78664 227773 78824 227807
rect 78664 227745 78699 227773
rect 78727 227745 78761 227773
rect 78789 227745 78824 227773
rect 78664 227728 78824 227745
rect 94024 227959 94184 227976
rect 94024 227931 94059 227959
rect 94087 227931 94121 227959
rect 94149 227931 94184 227959
rect 94024 227897 94184 227931
rect 94024 227869 94059 227897
rect 94087 227869 94121 227897
rect 94149 227869 94184 227897
rect 94024 227835 94184 227869
rect 94024 227807 94059 227835
rect 94087 227807 94121 227835
rect 94149 227807 94184 227835
rect 94024 227773 94184 227807
rect 94024 227745 94059 227773
rect 94087 227745 94121 227773
rect 94149 227745 94184 227773
rect 94024 227728 94184 227745
rect 109384 227959 109544 227976
rect 109384 227931 109419 227959
rect 109447 227931 109481 227959
rect 109509 227931 109544 227959
rect 109384 227897 109544 227931
rect 109384 227869 109419 227897
rect 109447 227869 109481 227897
rect 109509 227869 109544 227897
rect 109384 227835 109544 227869
rect 109384 227807 109419 227835
rect 109447 227807 109481 227835
rect 109509 227807 109544 227835
rect 109384 227773 109544 227807
rect 109384 227745 109419 227773
rect 109447 227745 109481 227773
rect 109509 227745 109544 227773
rect 109384 227728 109544 227745
rect 124744 227959 124904 227976
rect 124744 227931 124779 227959
rect 124807 227931 124841 227959
rect 124869 227931 124904 227959
rect 124744 227897 124904 227931
rect 124744 227869 124779 227897
rect 124807 227869 124841 227897
rect 124869 227869 124904 227897
rect 124744 227835 124904 227869
rect 124744 227807 124779 227835
rect 124807 227807 124841 227835
rect 124869 227807 124904 227835
rect 124744 227773 124904 227807
rect 124744 227745 124779 227773
rect 124807 227745 124841 227773
rect 124869 227745 124904 227773
rect 124744 227728 124904 227745
rect 140104 227959 140264 227976
rect 140104 227931 140139 227959
rect 140167 227931 140201 227959
rect 140229 227931 140264 227959
rect 140104 227897 140264 227931
rect 140104 227869 140139 227897
rect 140167 227869 140201 227897
rect 140229 227869 140264 227897
rect 140104 227835 140264 227869
rect 140104 227807 140139 227835
rect 140167 227807 140201 227835
rect 140229 227807 140264 227835
rect 140104 227773 140264 227807
rect 140104 227745 140139 227773
rect 140167 227745 140201 227773
rect 140229 227745 140264 227773
rect 140104 227728 140264 227745
rect 155464 227959 155624 227976
rect 155464 227931 155499 227959
rect 155527 227931 155561 227959
rect 155589 227931 155624 227959
rect 155464 227897 155624 227931
rect 155464 227869 155499 227897
rect 155527 227869 155561 227897
rect 155589 227869 155624 227897
rect 155464 227835 155624 227869
rect 155464 227807 155499 227835
rect 155527 227807 155561 227835
rect 155589 227807 155624 227835
rect 155464 227773 155624 227807
rect 155464 227745 155499 227773
rect 155527 227745 155561 227773
rect 155589 227745 155624 227773
rect 155464 227728 155624 227745
rect 170824 227959 170984 227976
rect 170824 227931 170859 227959
rect 170887 227931 170921 227959
rect 170949 227931 170984 227959
rect 170824 227897 170984 227931
rect 170824 227869 170859 227897
rect 170887 227869 170921 227897
rect 170949 227869 170984 227897
rect 170824 227835 170984 227869
rect 170824 227807 170859 227835
rect 170887 227807 170921 227835
rect 170949 227807 170984 227835
rect 170824 227773 170984 227807
rect 170824 227745 170859 227773
rect 170887 227745 170921 227773
rect 170949 227745 170984 227773
rect 170824 227728 170984 227745
rect 186184 227959 186344 227976
rect 186184 227931 186219 227959
rect 186247 227931 186281 227959
rect 186309 227931 186344 227959
rect 186184 227897 186344 227931
rect 186184 227869 186219 227897
rect 186247 227869 186281 227897
rect 186309 227869 186344 227897
rect 186184 227835 186344 227869
rect 186184 227807 186219 227835
rect 186247 227807 186281 227835
rect 186309 227807 186344 227835
rect 186184 227773 186344 227807
rect 186184 227745 186219 227773
rect 186247 227745 186281 227773
rect 186309 227745 186344 227773
rect 186184 227728 186344 227745
rect 201544 227959 201704 227976
rect 201544 227931 201579 227959
rect 201607 227931 201641 227959
rect 201669 227931 201704 227959
rect 201544 227897 201704 227931
rect 201544 227869 201579 227897
rect 201607 227869 201641 227897
rect 201669 227869 201704 227897
rect 201544 227835 201704 227869
rect 201544 227807 201579 227835
rect 201607 227807 201641 227835
rect 201669 227807 201704 227835
rect 201544 227773 201704 227807
rect 201544 227745 201579 227773
rect 201607 227745 201641 227773
rect 201669 227745 201704 227773
rect 201544 227728 201704 227745
rect 216904 227959 217064 227976
rect 216904 227931 216939 227959
rect 216967 227931 217001 227959
rect 217029 227931 217064 227959
rect 216904 227897 217064 227931
rect 216904 227869 216939 227897
rect 216967 227869 217001 227897
rect 217029 227869 217064 227897
rect 216904 227835 217064 227869
rect 216904 227807 216939 227835
rect 216967 227807 217001 227835
rect 217029 227807 217064 227835
rect 216904 227773 217064 227807
rect 216904 227745 216939 227773
rect 216967 227745 217001 227773
rect 217029 227745 217064 227773
rect 216904 227728 217064 227745
rect 232264 227959 232424 227976
rect 232264 227931 232299 227959
rect 232327 227931 232361 227959
rect 232389 227931 232424 227959
rect 232264 227897 232424 227931
rect 232264 227869 232299 227897
rect 232327 227869 232361 227897
rect 232389 227869 232424 227897
rect 232264 227835 232424 227869
rect 232264 227807 232299 227835
rect 232327 227807 232361 227835
rect 232389 227807 232424 227835
rect 232264 227773 232424 227807
rect 232264 227745 232299 227773
rect 232327 227745 232361 227773
rect 232389 227745 232424 227773
rect 232264 227728 232424 227745
rect 247624 227959 247784 227976
rect 247624 227931 247659 227959
rect 247687 227931 247721 227959
rect 247749 227931 247784 227959
rect 247624 227897 247784 227931
rect 247624 227869 247659 227897
rect 247687 227869 247721 227897
rect 247749 227869 247784 227897
rect 247624 227835 247784 227869
rect 247624 227807 247659 227835
rect 247687 227807 247721 227835
rect 247749 227807 247784 227835
rect 247624 227773 247784 227807
rect 247624 227745 247659 227773
rect 247687 227745 247721 227773
rect 247749 227745 247784 227773
rect 247624 227728 247784 227745
rect 254529 227959 254839 236745
rect 254529 227931 254577 227959
rect 254605 227931 254639 227959
rect 254667 227931 254701 227959
rect 254729 227931 254763 227959
rect 254791 227931 254839 227959
rect 254529 227897 254839 227931
rect 254529 227869 254577 227897
rect 254605 227869 254639 227897
rect 254667 227869 254701 227897
rect 254729 227869 254763 227897
rect 254791 227869 254839 227897
rect 254529 227835 254839 227869
rect 254529 227807 254577 227835
rect 254605 227807 254639 227835
rect 254667 227807 254701 227835
rect 254729 227807 254763 227835
rect 254791 227807 254839 227835
rect 254529 227773 254839 227807
rect 254529 227745 254577 227773
rect 254605 227745 254639 227773
rect 254667 227745 254701 227773
rect 254729 227745 254763 227773
rect 254791 227745 254839 227773
rect 31389 221931 31437 221959
rect 31465 221931 31499 221959
rect 31527 221931 31561 221959
rect 31589 221931 31623 221959
rect 31651 221931 31699 221959
rect 31389 221897 31699 221931
rect 31389 221869 31437 221897
rect 31465 221869 31499 221897
rect 31527 221869 31561 221897
rect 31589 221869 31623 221897
rect 31651 221869 31699 221897
rect 31389 221835 31699 221869
rect 31389 221807 31437 221835
rect 31465 221807 31499 221835
rect 31527 221807 31561 221835
rect 31589 221807 31623 221835
rect 31651 221807 31699 221835
rect 31389 221773 31699 221807
rect 31389 221745 31437 221773
rect 31465 221745 31499 221773
rect 31527 221745 31561 221773
rect 31589 221745 31623 221773
rect 31651 221745 31699 221773
rect 31389 212959 31699 221745
rect 40264 221959 40424 221976
rect 40264 221931 40299 221959
rect 40327 221931 40361 221959
rect 40389 221931 40424 221959
rect 40264 221897 40424 221931
rect 40264 221869 40299 221897
rect 40327 221869 40361 221897
rect 40389 221869 40424 221897
rect 40264 221835 40424 221869
rect 40264 221807 40299 221835
rect 40327 221807 40361 221835
rect 40389 221807 40424 221835
rect 40264 221773 40424 221807
rect 40264 221745 40299 221773
rect 40327 221745 40361 221773
rect 40389 221745 40424 221773
rect 40264 221728 40424 221745
rect 55624 221959 55784 221976
rect 55624 221931 55659 221959
rect 55687 221931 55721 221959
rect 55749 221931 55784 221959
rect 55624 221897 55784 221931
rect 55624 221869 55659 221897
rect 55687 221869 55721 221897
rect 55749 221869 55784 221897
rect 55624 221835 55784 221869
rect 55624 221807 55659 221835
rect 55687 221807 55721 221835
rect 55749 221807 55784 221835
rect 55624 221773 55784 221807
rect 55624 221745 55659 221773
rect 55687 221745 55721 221773
rect 55749 221745 55784 221773
rect 55624 221728 55784 221745
rect 70984 221959 71144 221976
rect 70984 221931 71019 221959
rect 71047 221931 71081 221959
rect 71109 221931 71144 221959
rect 70984 221897 71144 221931
rect 70984 221869 71019 221897
rect 71047 221869 71081 221897
rect 71109 221869 71144 221897
rect 70984 221835 71144 221869
rect 70984 221807 71019 221835
rect 71047 221807 71081 221835
rect 71109 221807 71144 221835
rect 70984 221773 71144 221807
rect 70984 221745 71019 221773
rect 71047 221745 71081 221773
rect 71109 221745 71144 221773
rect 70984 221728 71144 221745
rect 86344 221959 86504 221976
rect 86344 221931 86379 221959
rect 86407 221931 86441 221959
rect 86469 221931 86504 221959
rect 86344 221897 86504 221931
rect 86344 221869 86379 221897
rect 86407 221869 86441 221897
rect 86469 221869 86504 221897
rect 86344 221835 86504 221869
rect 86344 221807 86379 221835
rect 86407 221807 86441 221835
rect 86469 221807 86504 221835
rect 86344 221773 86504 221807
rect 86344 221745 86379 221773
rect 86407 221745 86441 221773
rect 86469 221745 86504 221773
rect 86344 221728 86504 221745
rect 101704 221959 101864 221976
rect 101704 221931 101739 221959
rect 101767 221931 101801 221959
rect 101829 221931 101864 221959
rect 101704 221897 101864 221931
rect 101704 221869 101739 221897
rect 101767 221869 101801 221897
rect 101829 221869 101864 221897
rect 101704 221835 101864 221869
rect 101704 221807 101739 221835
rect 101767 221807 101801 221835
rect 101829 221807 101864 221835
rect 101704 221773 101864 221807
rect 101704 221745 101739 221773
rect 101767 221745 101801 221773
rect 101829 221745 101864 221773
rect 101704 221728 101864 221745
rect 117064 221959 117224 221976
rect 117064 221931 117099 221959
rect 117127 221931 117161 221959
rect 117189 221931 117224 221959
rect 117064 221897 117224 221931
rect 117064 221869 117099 221897
rect 117127 221869 117161 221897
rect 117189 221869 117224 221897
rect 117064 221835 117224 221869
rect 117064 221807 117099 221835
rect 117127 221807 117161 221835
rect 117189 221807 117224 221835
rect 117064 221773 117224 221807
rect 117064 221745 117099 221773
rect 117127 221745 117161 221773
rect 117189 221745 117224 221773
rect 117064 221728 117224 221745
rect 132424 221959 132584 221976
rect 132424 221931 132459 221959
rect 132487 221931 132521 221959
rect 132549 221931 132584 221959
rect 132424 221897 132584 221931
rect 132424 221869 132459 221897
rect 132487 221869 132521 221897
rect 132549 221869 132584 221897
rect 132424 221835 132584 221869
rect 132424 221807 132459 221835
rect 132487 221807 132521 221835
rect 132549 221807 132584 221835
rect 132424 221773 132584 221807
rect 132424 221745 132459 221773
rect 132487 221745 132521 221773
rect 132549 221745 132584 221773
rect 132424 221728 132584 221745
rect 147784 221959 147944 221976
rect 147784 221931 147819 221959
rect 147847 221931 147881 221959
rect 147909 221931 147944 221959
rect 147784 221897 147944 221931
rect 147784 221869 147819 221897
rect 147847 221869 147881 221897
rect 147909 221869 147944 221897
rect 147784 221835 147944 221869
rect 147784 221807 147819 221835
rect 147847 221807 147881 221835
rect 147909 221807 147944 221835
rect 147784 221773 147944 221807
rect 147784 221745 147819 221773
rect 147847 221745 147881 221773
rect 147909 221745 147944 221773
rect 147784 221728 147944 221745
rect 163144 221959 163304 221976
rect 163144 221931 163179 221959
rect 163207 221931 163241 221959
rect 163269 221931 163304 221959
rect 163144 221897 163304 221931
rect 163144 221869 163179 221897
rect 163207 221869 163241 221897
rect 163269 221869 163304 221897
rect 163144 221835 163304 221869
rect 163144 221807 163179 221835
rect 163207 221807 163241 221835
rect 163269 221807 163304 221835
rect 163144 221773 163304 221807
rect 163144 221745 163179 221773
rect 163207 221745 163241 221773
rect 163269 221745 163304 221773
rect 163144 221728 163304 221745
rect 178504 221959 178664 221976
rect 178504 221931 178539 221959
rect 178567 221931 178601 221959
rect 178629 221931 178664 221959
rect 178504 221897 178664 221931
rect 178504 221869 178539 221897
rect 178567 221869 178601 221897
rect 178629 221869 178664 221897
rect 178504 221835 178664 221869
rect 178504 221807 178539 221835
rect 178567 221807 178601 221835
rect 178629 221807 178664 221835
rect 178504 221773 178664 221807
rect 178504 221745 178539 221773
rect 178567 221745 178601 221773
rect 178629 221745 178664 221773
rect 178504 221728 178664 221745
rect 193864 221959 194024 221976
rect 193864 221931 193899 221959
rect 193927 221931 193961 221959
rect 193989 221931 194024 221959
rect 193864 221897 194024 221931
rect 193864 221869 193899 221897
rect 193927 221869 193961 221897
rect 193989 221869 194024 221897
rect 193864 221835 194024 221869
rect 193864 221807 193899 221835
rect 193927 221807 193961 221835
rect 193989 221807 194024 221835
rect 193864 221773 194024 221807
rect 193864 221745 193899 221773
rect 193927 221745 193961 221773
rect 193989 221745 194024 221773
rect 193864 221728 194024 221745
rect 209224 221959 209384 221976
rect 209224 221931 209259 221959
rect 209287 221931 209321 221959
rect 209349 221931 209384 221959
rect 209224 221897 209384 221931
rect 209224 221869 209259 221897
rect 209287 221869 209321 221897
rect 209349 221869 209384 221897
rect 209224 221835 209384 221869
rect 209224 221807 209259 221835
rect 209287 221807 209321 221835
rect 209349 221807 209384 221835
rect 209224 221773 209384 221807
rect 209224 221745 209259 221773
rect 209287 221745 209321 221773
rect 209349 221745 209384 221773
rect 209224 221728 209384 221745
rect 224584 221959 224744 221976
rect 224584 221931 224619 221959
rect 224647 221931 224681 221959
rect 224709 221931 224744 221959
rect 224584 221897 224744 221931
rect 224584 221869 224619 221897
rect 224647 221869 224681 221897
rect 224709 221869 224744 221897
rect 224584 221835 224744 221869
rect 224584 221807 224619 221835
rect 224647 221807 224681 221835
rect 224709 221807 224744 221835
rect 224584 221773 224744 221807
rect 224584 221745 224619 221773
rect 224647 221745 224681 221773
rect 224709 221745 224744 221773
rect 224584 221728 224744 221745
rect 239944 221959 240104 221976
rect 239944 221931 239979 221959
rect 240007 221931 240041 221959
rect 240069 221931 240104 221959
rect 239944 221897 240104 221931
rect 239944 221869 239979 221897
rect 240007 221869 240041 221897
rect 240069 221869 240104 221897
rect 239944 221835 240104 221869
rect 239944 221807 239979 221835
rect 240007 221807 240041 221835
rect 240069 221807 240104 221835
rect 239944 221773 240104 221807
rect 239944 221745 239979 221773
rect 240007 221745 240041 221773
rect 240069 221745 240104 221773
rect 239944 221728 240104 221745
rect 32584 218959 32744 218976
rect 32584 218931 32619 218959
rect 32647 218931 32681 218959
rect 32709 218931 32744 218959
rect 32584 218897 32744 218931
rect 32584 218869 32619 218897
rect 32647 218869 32681 218897
rect 32709 218869 32744 218897
rect 32584 218835 32744 218869
rect 32584 218807 32619 218835
rect 32647 218807 32681 218835
rect 32709 218807 32744 218835
rect 32584 218773 32744 218807
rect 32584 218745 32619 218773
rect 32647 218745 32681 218773
rect 32709 218745 32744 218773
rect 32584 218728 32744 218745
rect 47944 218959 48104 218976
rect 47944 218931 47979 218959
rect 48007 218931 48041 218959
rect 48069 218931 48104 218959
rect 47944 218897 48104 218931
rect 47944 218869 47979 218897
rect 48007 218869 48041 218897
rect 48069 218869 48104 218897
rect 47944 218835 48104 218869
rect 47944 218807 47979 218835
rect 48007 218807 48041 218835
rect 48069 218807 48104 218835
rect 47944 218773 48104 218807
rect 47944 218745 47979 218773
rect 48007 218745 48041 218773
rect 48069 218745 48104 218773
rect 47944 218728 48104 218745
rect 63304 218959 63464 218976
rect 63304 218931 63339 218959
rect 63367 218931 63401 218959
rect 63429 218931 63464 218959
rect 63304 218897 63464 218931
rect 63304 218869 63339 218897
rect 63367 218869 63401 218897
rect 63429 218869 63464 218897
rect 63304 218835 63464 218869
rect 63304 218807 63339 218835
rect 63367 218807 63401 218835
rect 63429 218807 63464 218835
rect 63304 218773 63464 218807
rect 63304 218745 63339 218773
rect 63367 218745 63401 218773
rect 63429 218745 63464 218773
rect 63304 218728 63464 218745
rect 78664 218959 78824 218976
rect 78664 218931 78699 218959
rect 78727 218931 78761 218959
rect 78789 218931 78824 218959
rect 78664 218897 78824 218931
rect 78664 218869 78699 218897
rect 78727 218869 78761 218897
rect 78789 218869 78824 218897
rect 78664 218835 78824 218869
rect 78664 218807 78699 218835
rect 78727 218807 78761 218835
rect 78789 218807 78824 218835
rect 78664 218773 78824 218807
rect 78664 218745 78699 218773
rect 78727 218745 78761 218773
rect 78789 218745 78824 218773
rect 78664 218728 78824 218745
rect 94024 218959 94184 218976
rect 94024 218931 94059 218959
rect 94087 218931 94121 218959
rect 94149 218931 94184 218959
rect 94024 218897 94184 218931
rect 94024 218869 94059 218897
rect 94087 218869 94121 218897
rect 94149 218869 94184 218897
rect 94024 218835 94184 218869
rect 94024 218807 94059 218835
rect 94087 218807 94121 218835
rect 94149 218807 94184 218835
rect 94024 218773 94184 218807
rect 94024 218745 94059 218773
rect 94087 218745 94121 218773
rect 94149 218745 94184 218773
rect 94024 218728 94184 218745
rect 109384 218959 109544 218976
rect 109384 218931 109419 218959
rect 109447 218931 109481 218959
rect 109509 218931 109544 218959
rect 109384 218897 109544 218931
rect 109384 218869 109419 218897
rect 109447 218869 109481 218897
rect 109509 218869 109544 218897
rect 109384 218835 109544 218869
rect 109384 218807 109419 218835
rect 109447 218807 109481 218835
rect 109509 218807 109544 218835
rect 109384 218773 109544 218807
rect 109384 218745 109419 218773
rect 109447 218745 109481 218773
rect 109509 218745 109544 218773
rect 109384 218728 109544 218745
rect 124744 218959 124904 218976
rect 124744 218931 124779 218959
rect 124807 218931 124841 218959
rect 124869 218931 124904 218959
rect 124744 218897 124904 218931
rect 124744 218869 124779 218897
rect 124807 218869 124841 218897
rect 124869 218869 124904 218897
rect 124744 218835 124904 218869
rect 124744 218807 124779 218835
rect 124807 218807 124841 218835
rect 124869 218807 124904 218835
rect 124744 218773 124904 218807
rect 124744 218745 124779 218773
rect 124807 218745 124841 218773
rect 124869 218745 124904 218773
rect 124744 218728 124904 218745
rect 140104 218959 140264 218976
rect 140104 218931 140139 218959
rect 140167 218931 140201 218959
rect 140229 218931 140264 218959
rect 140104 218897 140264 218931
rect 140104 218869 140139 218897
rect 140167 218869 140201 218897
rect 140229 218869 140264 218897
rect 140104 218835 140264 218869
rect 140104 218807 140139 218835
rect 140167 218807 140201 218835
rect 140229 218807 140264 218835
rect 140104 218773 140264 218807
rect 140104 218745 140139 218773
rect 140167 218745 140201 218773
rect 140229 218745 140264 218773
rect 140104 218728 140264 218745
rect 155464 218959 155624 218976
rect 155464 218931 155499 218959
rect 155527 218931 155561 218959
rect 155589 218931 155624 218959
rect 155464 218897 155624 218931
rect 155464 218869 155499 218897
rect 155527 218869 155561 218897
rect 155589 218869 155624 218897
rect 155464 218835 155624 218869
rect 155464 218807 155499 218835
rect 155527 218807 155561 218835
rect 155589 218807 155624 218835
rect 155464 218773 155624 218807
rect 155464 218745 155499 218773
rect 155527 218745 155561 218773
rect 155589 218745 155624 218773
rect 155464 218728 155624 218745
rect 170824 218959 170984 218976
rect 170824 218931 170859 218959
rect 170887 218931 170921 218959
rect 170949 218931 170984 218959
rect 170824 218897 170984 218931
rect 170824 218869 170859 218897
rect 170887 218869 170921 218897
rect 170949 218869 170984 218897
rect 170824 218835 170984 218869
rect 170824 218807 170859 218835
rect 170887 218807 170921 218835
rect 170949 218807 170984 218835
rect 170824 218773 170984 218807
rect 170824 218745 170859 218773
rect 170887 218745 170921 218773
rect 170949 218745 170984 218773
rect 170824 218728 170984 218745
rect 186184 218959 186344 218976
rect 186184 218931 186219 218959
rect 186247 218931 186281 218959
rect 186309 218931 186344 218959
rect 186184 218897 186344 218931
rect 186184 218869 186219 218897
rect 186247 218869 186281 218897
rect 186309 218869 186344 218897
rect 186184 218835 186344 218869
rect 186184 218807 186219 218835
rect 186247 218807 186281 218835
rect 186309 218807 186344 218835
rect 186184 218773 186344 218807
rect 186184 218745 186219 218773
rect 186247 218745 186281 218773
rect 186309 218745 186344 218773
rect 186184 218728 186344 218745
rect 201544 218959 201704 218976
rect 201544 218931 201579 218959
rect 201607 218931 201641 218959
rect 201669 218931 201704 218959
rect 201544 218897 201704 218931
rect 201544 218869 201579 218897
rect 201607 218869 201641 218897
rect 201669 218869 201704 218897
rect 201544 218835 201704 218869
rect 201544 218807 201579 218835
rect 201607 218807 201641 218835
rect 201669 218807 201704 218835
rect 201544 218773 201704 218807
rect 201544 218745 201579 218773
rect 201607 218745 201641 218773
rect 201669 218745 201704 218773
rect 201544 218728 201704 218745
rect 216904 218959 217064 218976
rect 216904 218931 216939 218959
rect 216967 218931 217001 218959
rect 217029 218931 217064 218959
rect 216904 218897 217064 218931
rect 216904 218869 216939 218897
rect 216967 218869 217001 218897
rect 217029 218869 217064 218897
rect 216904 218835 217064 218869
rect 216904 218807 216939 218835
rect 216967 218807 217001 218835
rect 217029 218807 217064 218835
rect 216904 218773 217064 218807
rect 216904 218745 216939 218773
rect 216967 218745 217001 218773
rect 217029 218745 217064 218773
rect 216904 218728 217064 218745
rect 232264 218959 232424 218976
rect 232264 218931 232299 218959
rect 232327 218931 232361 218959
rect 232389 218931 232424 218959
rect 232264 218897 232424 218931
rect 232264 218869 232299 218897
rect 232327 218869 232361 218897
rect 232389 218869 232424 218897
rect 232264 218835 232424 218869
rect 232264 218807 232299 218835
rect 232327 218807 232361 218835
rect 232389 218807 232424 218835
rect 232264 218773 232424 218807
rect 232264 218745 232299 218773
rect 232327 218745 232361 218773
rect 232389 218745 232424 218773
rect 232264 218728 232424 218745
rect 247624 218959 247784 218976
rect 247624 218931 247659 218959
rect 247687 218931 247721 218959
rect 247749 218931 247784 218959
rect 247624 218897 247784 218931
rect 247624 218869 247659 218897
rect 247687 218869 247721 218897
rect 247749 218869 247784 218897
rect 247624 218835 247784 218869
rect 247624 218807 247659 218835
rect 247687 218807 247721 218835
rect 247749 218807 247784 218835
rect 247624 218773 247784 218807
rect 247624 218745 247659 218773
rect 247687 218745 247721 218773
rect 247749 218745 247784 218773
rect 247624 218728 247784 218745
rect 254529 218959 254839 227745
rect 254529 218931 254577 218959
rect 254605 218931 254639 218959
rect 254667 218931 254701 218959
rect 254729 218931 254763 218959
rect 254791 218931 254839 218959
rect 254529 218897 254839 218931
rect 254529 218869 254577 218897
rect 254605 218869 254639 218897
rect 254667 218869 254701 218897
rect 254729 218869 254763 218897
rect 254791 218869 254839 218897
rect 254529 218835 254839 218869
rect 254529 218807 254577 218835
rect 254605 218807 254639 218835
rect 254667 218807 254701 218835
rect 254729 218807 254763 218835
rect 254791 218807 254839 218835
rect 254529 218773 254839 218807
rect 254529 218745 254577 218773
rect 254605 218745 254639 218773
rect 254667 218745 254701 218773
rect 254729 218745 254763 218773
rect 254791 218745 254839 218773
rect 31389 212931 31437 212959
rect 31465 212931 31499 212959
rect 31527 212931 31561 212959
rect 31589 212931 31623 212959
rect 31651 212931 31699 212959
rect 31389 212897 31699 212931
rect 31389 212869 31437 212897
rect 31465 212869 31499 212897
rect 31527 212869 31561 212897
rect 31589 212869 31623 212897
rect 31651 212869 31699 212897
rect 31389 212835 31699 212869
rect 31389 212807 31437 212835
rect 31465 212807 31499 212835
rect 31527 212807 31561 212835
rect 31589 212807 31623 212835
rect 31651 212807 31699 212835
rect 31389 212773 31699 212807
rect 31389 212745 31437 212773
rect 31465 212745 31499 212773
rect 31527 212745 31561 212773
rect 31589 212745 31623 212773
rect 31651 212745 31699 212773
rect 31389 203959 31699 212745
rect 40264 212959 40424 212976
rect 40264 212931 40299 212959
rect 40327 212931 40361 212959
rect 40389 212931 40424 212959
rect 40264 212897 40424 212931
rect 40264 212869 40299 212897
rect 40327 212869 40361 212897
rect 40389 212869 40424 212897
rect 40264 212835 40424 212869
rect 40264 212807 40299 212835
rect 40327 212807 40361 212835
rect 40389 212807 40424 212835
rect 40264 212773 40424 212807
rect 40264 212745 40299 212773
rect 40327 212745 40361 212773
rect 40389 212745 40424 212773
rect 40264 212728 40424 212745
rect 55624 212959 55784 212976
rect 55624 212931 55659 212959
rect 55687 212931 55721 212959
rect 55749 212931 55784 212959
rect 55624 212897 55784 212931
rect 55624 212869 55659 212897
rect 55687 212869 55721 212897
rect 55749 212869 55784 212897
rect 55624 212835 55784 212869
rect 55624 212807 55659 212835
rect 55687 212807 55721 212835
rect 55749 212807 55784 212835
rect 55624 212773 55784 212807
rect 55624 212745 55659 212773
rect 55687 212745 55721 212773
rect 55749 212745 55784 212773
rect 55624 212728 55784 212745
rect 70984 212959 71144 212976
rect 70984 212931 71019 212959
rect 71047 212931 71081 212959
rect 71109 212931 71144 212959
rect 70984 212897 71144 212931
rect 70984 212869 71019 212897
rect 71047 212869 71081 212897
rect 71109 212869 71144 212897
rect 70984 212835 71144 212869
rect 70984 212807 71019 212835
rect 71047 212807 71081 212835
rect 71109 212807 71144 212835
rect 70984 212773 71144 212807
rect 70984 212745 71019 212773
rect 71047 212745 71081 212773
rect 71109 212745 71144 212773
rect 70984 212728 71144 212745
rect 86344 212959 86504 212976
rect 86344 212931 86379 212959
rect 86407 212931 86441 212959
rect 86469 212931 86504 212959
rect 86344 212897 86504 212931
rect 86344 212869 86379 212897
rect 86407 212869 86441 212897
rect 86469 212869 86504 212897
rect 86344 212835 86504 212869
rect 86344 212807 86379 212835
rect 86407 212807 86441 212835
rect 86469 212807 86504 212835
rect 86344 212773 86504 212807
rect 86344 212745 86379 212773
rect 86407 212745 86441 212773
rect 86469 212745 86504 212773
rect 86344 212728 86504 212745
rect 101704 212959 101864 212976
rect 101704 212931 101739 212959
rect 101767 212931 101801 212959
rect 101829 212931 101864 212959
rect 101704 212897 101864 212931
rect 101704 212869 101739 212897
rect 101767 212869 101801 212897
rect 101829 212869 101864 212897
rect 101704 212835 101864 212869
rect 101704 212807 101739 212835
rect 101767 212807 101801 212835
rect 101829 212807 101864 212835
rect 101704 212773 101864 212807
rect 101704 212745 101739 212773
rect 101767 212745 101801 212773
rect 101829 212745 101864 212773
rect 101704 212728 101864 212745
rect 117064 212959 117224 212976
rect 117064 212931 117099 212959
rect 117127 212931 117161 212959
rect 117189 212931 117224 212959
rect 117064 212897 117224 212931
rect 117064 212869 117099 212897
rect 117127 212869 117161 212897
rect 117189 212869 117224 212897
rect 117064 212835 117224 212869
rect 117064 212807 117099 212835
rect 117127 212807 117161 212835
rect 117189 212807 117224 212835
rect 117064 212773 117224 212807
rect 117064 212745 117099 212773
rect 117127 212745 117161 212773
rect 117189 212745 117224 212773
rect 117064 212728 117224 212745
rect 132424 212959 132584 212976
rect 132424 212931 132459 212959
rect 132487 212931 132521 212959
rect 132549 212931 132584 212959
rect 132424 212897 132584 212931
rect 132424 212869 132459 212897
rect 132487 212869 132521 212897
rect 132549 212869 132584 212897
rect 132424 212835 132584 212869
rect 132424 212807 132459 212835
rect 132487 212807 132521 212835
rect 132549 212807 132584 212835
rect 132424 212773 132584 212807
rect 132424 212745 132459 212773
rect 132487 212745 132521 212773
rect 132549 212745 132584 212773
rect 132424 212728 132584 212745
rect 147784 212959 147944 212976
rect 147784 212931 147819 212959
rect 147847 212931 147881 212959
rect 147909 212931 147944 212959
rect 147784 212897 147944 212931
rect 147784 212869 147819 212897
rect 147847 212869 147881 212897
rect 147909 212869 147944 212897
rect 147784 212835 147944 212869
rect 147784 212807 147819 212835
rect 147847 212807 147881 212835
rect 147909 212807 147944 212835
rect 147784 212773 147944 212807
rect 147784 212745 147819 212773
rect 147847 212745 147881 212773
rect 147909 212745 147944 212773
rect 147784 212728 147944 212745
rect 163144 212959 163304 212976
rect 163144 212931 163179 212959
rect 163207 212931 163241 212959
rect 163269 212931 163304 212959
rect 163144 212897 163304 212931
rect 163144 212869 163179 212897
rect 163207 212869 163241 212897
rect 163269 212869 163304 212897
rect 163144 212835 163304 212869
rect 163144 212807 163179 212835
rect 163207 212807 163241 212835
rect 163269 212807 163304 212835
rect 163144 212773 163304 212807
rect 163144 212745 163179 212773
rect 163207 212745 163241 212773
rect 163269 212745 163304 212773
rect 163144 212728 163304 212745
rect 178504 212959 178664 212976
rect 178504 212931 178539 212959
rect 178567 212931 178601 212959
rect 178629 212931 178664 212959
rect 178504 212897 178664 212931
rect 178504 212869 178539 212897
rect 178567 212869 178601 212897
rect 178629 212869 178664 212897
rect 178504 212835 178664 212869
rect 178504 212807 178539 212835
rect 178567 212807 178601 212835
rect 178629 212807 178664 212835
rect 178504 212773 178664 212807
rect 178504 212745 178539 212773
rect 178567 212745 178601 212773
rect 178629 212745 178664 212773
rect 178504 212728 178664 212745
rect 193864 212959 194024 212976
rect 193864 212931 193899 212959
rect 193927 212931 193961 212959
rect 193989 212931 194024 212959
rect 193864 212897 194024 212931
rect 193864 212869 193899 212897
rect 193927 212869 193961 212897
rect 193989 212869 194024 212897
rect 193864 212835 194024 212869
rect 193864 212807 193899 212835
rect 193927 212807 193961 212835
rect 193989 212807 194024 212835
rect 193864 212773 194024 212807
rect 193864 212745 193899 212773
rect 193927 212745 193961 212773
rect 193989 212745 194024 212773
rect 193864 212728 194024 212745
rect 209224 212959 209384 212976
rect 209224 212931 209259 212959
rect 209287 212931 209321 212959
rect 209349 212931 209384 212959
rect 209224 212897 209384 212931
rect 209224 212869 209259 212897
rect 209287 212869 209321 212897
rect 209349 212869 209384 212897
rect 209224 212835 209384 212869
rect 209224 212807 209259 212835
rect 209287 212807 209321 212835
rect 209349 212807 209384 212835
rect 209224 212773 209384 212807
rect 209224 212745 209259 212773
rect 209287 212745 209321 212773
rect 209349 212745 209384 212773
rect 209224 212728 209384 212745
rect 224584 212959 224744 212976
rect 224584 212931 224619 212959
rect 224647 212931 224681 212959
rect 224709 212931 224744 212959
rect 224584 212897 224744 212931
rect 224584 212869 224619 212897
rect 224647 212869 224681 212897
rect 224709 212869 224744 212897
rect 224584 212835 224744 212869
rect 224584 212807 224619 212835
rect 224647 212807 224681 212835
rect 224709 212807 224744 212835
rect 224584 212773 224744 212807
rect 224584 212745 224619 212773
rect 224647 212745 224681 212773
rect 224709 212745 224744 212773
rect 224584 212728 224744 212745
rect 239944 212959 240104 212976
rect 239944 212931 239979 212959
rect 240007 212931 240041 212959
rect 240069 212931 240104 212959
rect 239944 212897 240104 212931
rect 239944 212869 239979 212897
rect 240007 212869 240041 212897
rect 240069 212869 240104 212897
rect 239944 212835 240104 212869
rect 239944 212807 239979 212835
rect 240007 212807 240041 212835
rect 240069 212807 240104 212835
rect 239944 212773 240104 212807
rect 239944 212745 239979 212773
rect 240007 212745 240041 212773
rect 240069 212745 240104 212773
rect 239944 212728 240104 212745
rect 32584 209959 32744 209976
rect 32584 209931 32619 209959
rect 32647 209931 32681 209959
rect 32709 209931 32744 209959
rect 32584 209897 32744 209931
rect 32584 209869 32619 209897
rect 32647 209869 32681 209897
rect 32709 209869 32744 209897
rect 32584 209835 32744 209869
rect 32584 209807 32619 209835
rect 32647 209807 32681 209835
rect 32709 209807 32744 209835
rect 32584 209773 32744 209807
rect 32584 209745 32619 209773
rect 32647 209745 32681 209773
rect 32709 209745 32744 209773
rect 32584 209728 32744 209745
rect 47944 209959 48104 209976
rect 47944 209931 47979 209959
rect 48007 209931 48041 209959
rect 48069 209931 48104 209959
rect 47944 209897 48104 209931
rect 47944 209869 47979 209897
rect 48007 209869 48041 209897
rect 48069 209869 48104 209897
rect 47944 209835 48104 209869
rect 47944 209807 47979 209835
rect 48007 209807 48041 209835
rect 48069 209807 48104 209835
rect 47944 209773 48104 209807
rect 47944 209745 47979 209773
rect 48007 209745 48041 209773
rect 48069 209745 48104 209773
rect 47944 209728 48104 209745
rect 63304 209959 63464 209976
rect 63304 209931 63339 209959
rect 63367 209931 63401 209959
rect 63429 209931 63464 209959
rect 63304 209897 63464 209931
rect 63304 209869 63339 209897
rect 63367 209869 63401 209897
rect 63429 209869 63464 209897
rect 63304 209835 63464 209869
rect 63304 209807 63339 209835
rect 63367 209807 63401 209835
rect 63429 209807 63464 209835
rect 63304 209773 63464 209807
rect 63304 209745 63339 209773
rect 63367 209745 63401 209773
rect 63429 209745 63464 209773
rect 63304 209728 63464 209745
rect 78664 209959 78824 209976
rect 78664 209931 78699 209959
rect 78727 209931 78761 209959
rect 78789 209931 78824 209959
rect 78664 209897 78824 209931
rect 78664 209869 78699 209897
rect 78727 209869 78761 209897
rect 78789 209869 78824 209897
rect 78664 209835 78824 209869
rect 78664 209807 78699 209835
rect 78727 209807 78761 209835
rect 78789 209807 78824 209835
rect 78664 209773 78824 209807
rect 78664 209745 78699 209773
rect 78727 209745 78761 209773
rect 78789 209745 78824 209773
rect 78664 209728 78824 209745
rect 94024 209959 94184 209976
rect 94024 209931 94059 209959
rect 94087 209931 94121 209959
rect 94149 209931 94184 209959
rect 94024 209897 94184 209931
rect 94024 209869 94059 209897
rect 94087 209869 94121 209897
rect 94149 209869 94184 209897
rect 94024 209835 94184 209869
rect 94024 209807 94059 209835
rect 94087 209807 94121 209835
rect 94149 209807 94184 209835
rect 94024 209773 94184 209807
rect 94024 209745 94059 209773
rect 94087 209745 94121 209773
rect 94149 209745 94184 209773
rect 94024 209728 94184 209745
rect 109384 209959 109544 209976
rect 109384 209931 109419 209959
rect 109447 209931 109481 209959
rect 109509 209931 109544 209959
rect 109384 209897 109544 209931
rect 109384 209869 109419 209897
rect 109447 209869 109481 209897
rect 109509 209869 109544 209897
rect 109384 209835 109544 209869
rect 109384 209807 109419 209835
rect 109447 209807 109481 209835
rect 109509 209807 109544 209835
rect 109384 209773 109544 209807
rect 109384 209745 109419 209773
rect 109447 209745 109481 209773
rect 109509 209745 109544 209773
rect 109384 209728 109544 209745
rect 124744 209959 124904 209976
rect 124744 209931 124779 209959
rect 124807 209931 124841 209959
rect 124869 209931 124904 209959
rect 124744 209897 124904 209931
rect 124744 209869 124779 209897
rect 124807 209869 124841 209897
rect 124869 209869 124904 209897
rect 124744 209835 124904 209869
rect 124744 209807 124779 209835
rect 124807 209807 124841 209835
rect 124869 209807 124904 209835
rect 124744 209773 124904 209807
rect 124744 209745 124779 209773
rect 124807 209745 124841 209773
rect 124869 209745 124904 209773
rect 124744 209728 124904 209745
rect 140104 209959 140264 209976
rect 140104 209931 140139 209959
rect 140167 209931 140201 209959
rect 140229 209931 140264 209959
rect 140104 209897 140264 209931
rect 140104 209869 140139 209897
rect 140167 209869 140201 209897
rect 140229 209869 140264 209897
rect 140104 209835 140264 209869
rect 140104 209807 140139 209835
rect 140167 209807 140201 209835
rect 140229 209807 140264 209835
rect 140104 209773 140264 209807
rect 140104 209745 140139 209773
rect 140167 209745 140201 209773
rect 140229 209745 140264 209773
rect 140104 209728 140264 209745
rect 155464 209959 155624 209976
rect 155464 209931 155499 209959
rect 155527 209931 155561 209959
rect 155589 209931 155624 209959
rect 155464 209897 155624 209931
rect 155464 209869 155499 209897
rect 155527 209869 155561 209897
rect 155589 209869 155624 209897
rect 155464 209835 155624 209869
rect 155464 209807 155499 209835
rect 155527 209807 155561 209835
rect 155589 209807 155624 209835
rect 155464 209773 155624 209807
rect 155464 209745 155499 209773
rect 155527 209745 155561 209773
rect 155589 209745 155624 209773
rect 155464 209728 155624 209745
rect 170824 209959 170984 209976
rect 170824 209931 170859 209959
rect 170887 209931 170921 209959
rect 170949 209931 170984 209959
rect 170824 209897 170984 209931
rect 170824 209869 170859 209897
rect 170887 209869 170921 209897
rect 170949 209869 170984 209897
rect 170824 209835 170984 209869
rect 170824 209807 170859 209835
rect 170887 209807 170921 209835
rect 170949 209807 170984 209835
rect 170824 209773 170984 209807
rect 170824 209745 170859 209773
rect 170887 209745 170921 209773
rect 170949 209745 170984 209773
rect 170824 209728 170984 209745
rect 186184 209959 186344 209976
rect 186184 209931 186219 209959
rect 186247 209931 186281 209959
rect 186309 209931 186344 209959
rect 186184 209897 186344 209931
rect 186184 209869 186219 209897
rect 186247 209869 186281 209897
rect 186309 209869 186344 209897
rect 186184 209835 186344 209869
rect 186184 209807 186219 209835
rect 186247 209807 186281 209835
rect 186309 209807 186344 209835
rect 186184 209773 186344 209807
rect 186184 209745 186219 209773
rect 186247 209745 186281 209773
rect 186309 209745 186344 209773
rect 186184 209728 186344 209745
rect 201544 209959 201704 209976
rect 201544 209931 201579 209959
rect 201607 209931 201641 209959
rect 201669 209931 201704 209959
rect 201544 209897 201704 209931
rect 201544 209869 201579 209897
rect 201607 209869 201641 209897
rect 201669 209869 201704 209897
rect 201544 209835 201704 209869
rect 201544 209807 201579 209835
rect 201607 209807 201641 209835
rect 201669 209807 201704 209835
rect 201544 209773 201704 209807
rect 201544 209745 201579 209773
rect 201607 209745 201641 209773
rect 201669 209745 201704 209773
rect 201544 209728 201704 209745
rect 216904 209959 217064 209976
rect 216904 209931 216939 209959
rect 216967 209931 217001 209959
rect 217029 209931 217064 209959
rect 216904 209897 217064 209931
rect 216904 209869 216939 209897
rect 216967 209869 217001 209897
rect 217029 209869 217064 209897
rect 216904 209835 217064 209869
rect 216904 209807 216939 209835
rect 216967 209807 217001 209835
rect 217029 209807 217064 209835
rect 216904 209773 217064 209807
rect 216904 209745 216939 209773
rect 216967 209745 217001 209773
rect 217029 209745 217064 209773
rect 216904 209728 217064 209745
rect 232264 209959 232424 209976
rect 232264 209931 232299 209959
rect 232327 209931 232361 209959
rect 232389 209931 232424 209959
rect 232264 209897 232424 209931
rect 232264 209869 232299 209897
rect 232327 209869 232361 209897
rect 232389 209869 232424 209897
rect 232264 209835 232424 209869
rect 232264 209807 232299 209835
rect 232327 209807 232361 209835
rect 232389 209807 232424 209835
rect 232264 209773 232424 209807
rect 232264 209745 232299 209773
rect 232327 209745 232361 209773
rect 232389 209745 232424 209773
rect 232264 209728 232424 209745
rect 247624 209959 247784 209976
rect 247624 209931 247659 209959
rect 247687 209931 247721 209959
rect 247749 209931 247784 209959
rect 247624 209897 247784 209931
rect 247624 209869 247659 209897
rect 247687 209869 247721 209897
rect 247749 209869 247784 209897
rect 247624 209835 247784 209869
rect 247624 209807 247659 209835
rect 247687 209807 247721 209835
rect 247749 209807 247784 209835
rect 247624 209773 247784 209807
rect 247624 209745 247659 209773
rect 247687 209745 247721 209773
rect 247749 209745 247784 209773
rect 247624 209728 247784 209745
rect 254529 209959 254839 218745
rect 254529 209931 254577 209959
rect 254605 209931 254639 209959
rect 254667 209931 254701 209959
rect 254729 209931 254763 209959
rect 254791 209931 254839 209959
rect 254529 209897 254839 209931
rect 254529 209869 254577 209897
rect 254605 209869 254639 209897
rect 254667 209869 254701 209897
rect 254729 209869 254763 209897
rect 254791 209869 254839 209897
rect 254529 209835 254839 209869
rect 254529 209807 254577 209835
rect 254605 209807 254639 209835
rect 254667 209807 254701 209835
rect 254729 209807 254763 209835
rect 254791 209807 254839 209835
rect 254529 209773 254839 209807
rect 254529 209745 254577 209773
rect 254605 209745 254639 209773
rect 254667 209745 254701 209773
rect 254729 209745 254763 209773
rect 254791 209745 254839 209773
rect 31389 203931 31437 203959
rect 31465 203931 31499 203959
rect 31527 203931 31561 203959
rect 31589 203931 31623 203959
rect 31651 203931 31699 203959
rect 31389 203897 31699 203931
rect 31389 203869 31437 203897
rect 31465 203869 31499 203897
rect 31527 203869 31561 203897
rect 31589 203869 31623 203897
rect 31651 203869 31699 203897
rect 31389 203835 31699 203869
rect 31389 203807 31437 203835
rect 31465 203807 31499 203835
rect 31527 203807 31561 203835
rect 31589 203807 31623 203835
rect 31651 203807 31699 203835
rect 31389 203773 31699 203807
rect 31389 203745 31437 203773
rect 31465 203745 31499 203773
rect 31527 203745 31561 203773
rect 31589 203745 31623 203773
rect 31651 203745 31699 203773
rect 31389 194959 31699 203745
rect 40264 203959 40424 203976
rect 40264 203931 40299 203959
rect 40327 203931 40361 203959
rect 40389 203931 40424 203959
rect 40264 203897 40424 203931
rect 40264 203869 40299 203897
rect 40327 203869 40361 203897
rect 40389 203869 40424 203897
rect 40264 203835 40424 203869
rect 40264 203807 40299 203835
rect 40327 203807 40361 203835
rect 40389 203807 40424 203835
rect 40264 203773 40424 203807
rect 40264 203745 40299 203773
rect 40327 203745 40361 203773
rect 40389 203745 40424 203773
rect 40264 203728 40424 203745
rect 55624 203959 55784 203976
rect 55624 203931 55659 203959
rect 55687 203931 55721 203959
rect 55749 203931 55784 203959
rect 55624 203897 55784 203931
rect 55624 203869 55659 203897
rect 55687 203869 55721 203897
rect 55749 203869 55784 203897
rect 55624 203835 55784 203869
rect 55624 203807 55659 203835
rect 55687 203807 55721 203835
rect 55749 203807 55784 203835
rect 55624 203773 55784 203807
rect 55624 203745 55659 203773
rect 55687 203745 55721 203773
rect 55749 203745 55784 203773
rect 55624 203728 55784 203745
rect 70984 203959 71144 203976
rect 70984 203931 71019 203959
rect 71047 203931 71081 203959
rect 71109 203931 71144 203959
rect 70984 203897 71144 203931
rect 70984 203869 71019 203897
rect 71047 203869 71081 203897
rect 71109 203869 71144 203897
rect 70984 203835 71144 203869
rect 70984 203807 71019 203835
rect 71047 203807 71081 203835
rect 71109 203807 71144 203835
rect 70984 203773 71144 203807
rect 70984 203745 71019 203773
rect 71047 203745 71081 203773
rect 71109 203745 71144 203773
rect 70984 203728 71144 203745
rect 86344 203959 86504 203976
rect 86344 203931 86379 203959
rect 86407 203931 86441 203959
rect 86469 203931 86504 203959
rect 86344 203897 86504 203931
rect 86344 203869 86379 203897
rect 86407 203869 86441 203897
rect 86469 203869 86504 203897
rect 86344 203835 86504 203869
rect 86344 203807 86379 203835
rect 86407 203807 86441 203835
rect 86469 203807 86504 203835
rect 86344 203773 86504 203807
rect 86344 203745 86379 203773
rect 86407 203745 86441 203773
rect 86469 203745 86504 203773
rect 86344 203728 86504 203745
rect 101704 203959 101864 203976
rect 101704 203931 101739 203959
rect 101767 203931 101801 203959
rect 101829 203931 101864 203959
rect 101704 203897 101864 203931
rect 101704 203869 101739 203897
rect 101767 203869 101801 203897
rect 101829 203869 101864 203897
rect 101704 203835 101864 203869
rect 101704 203807 101739 203835
rect 101767 203807 101801 203835
rect 101829 203807 101864 203835
rect 101704 203773 101864 203807
rect 101704 203745 101739 203773
rect 101767 203745 101801 203773
rect 101829 203745 101864 203773
rect 101704 203728 101864 203745
rect 117064 203959 117224 203976
rect 117064 203931 117099 203959
rect 117127 203931 117161 203959
rect 117189 203931 117224 203959
rect 117064 203897 117224 203931
rect 117064 203869 117099 203897
rect 117127 203869 117161 203897
rect 117189 203869 117224 203897
rect 117064 203835 117224 203869
rect 117064 203807 117099 203835
rect 117127 203807 117161 203835
rect 117189 203807 117224 203835
rect 117064 203773 117224 203807
rect 117064 203745 117099 203773
rect 117127 203745 117161 203773
rect 117189 203745 117224 203773
rect 117064 203728 117224 203745
rect 132424 203959 132584 203976
rect 132424 203931 132459 203959
rect 132487 203931 132521 203959
rect 132549 203931 132584 203959
rect 132424 203897 132584 203931
rect 132424 203869 132459 203897
rect 132487 203869 132521 203897
rect 132549 203869 132584 203897
rect 132424 203835 132584 203869
rect 132424 203807 132459 203835
rect 132487 203807 132521 203835
rect 132549 203807 132584 203835
rect 132424 203773 132584 203807
rect 132424 203745 132459 203773
rect 132487 203745 132521 203773
rect 132549 203745 132584 203773
rect 132424 203728 132584 203745
rect 147784 203959 147944 203976
rect 147784 203931 147819 203959
rect 147847 203931 147881 203959
rect 147909 203931 147944 203959
rect 147784 203897 147944 203931
rect 147784 203869 147819 203897
rect 147847 203869 147881 203897
rect 147909 203869 147944 203897
rect 147784 203835 147944 203869
rect 147784 203807 147819 203835
rect 147847 203807 147881 203835
rect 147909 203807 147944 203835
rect 147784 203773 147944 203807
rect 147784 203745 147819 203773
rect 147847 203745 147881 203773
rect 147909 203745 147944 203773
rect 147784 203728 147944 203745
rect 163144 203959 163304 203976
rect 163144 203931 163179 203959
rect 163207 203931 163241 203959
rect 163269 203931 163304 203959
rect 163144 203897 163304 203931
rect 163144 203869 163179 203897
rect 163207 203869 163241 203897
rect 163269 203869 163304 203897
rect 163144 203835 163304 203869
rect 163144 203807 163179 203835
rect 163207 203807 163241 203835
rect 163269 203807 163304 203835
rect 163144 203773 163304 203807
rect 163144 203745 163179 203773
rect 163207 203745 163241 203773
rect 163269 203745 163304 203773
rect 163144 203728 163304 203745
rect 178504 203959 178664 203976
rect 178504 203931 178539 203959
rect 178567 203931 178601 203959
rect 178629 203931 178664 203959
rect 178504 203897 178664 203931
rect 178504 203869 178539 203897
rect 178567 203869 178601 203897
rect 178629 203869 178664 203897
rect 178504 203835 178664 203869
rect 178504 203807 178539 203835
rect 178567 203807 178601 203835
rect 178629 203807 178664 203835
rect 178504 203773 178664 203807
rect 178504 203745 178539 203773
rect 178567 203745 178601 203773
rect 178629 203745 178664 203773
rect 178504 203728 178664 203745
rect 193864 203959 194024 203976
rect 193864 203931 193899 203959
rect 193927 203931 193961 203959
rect 193989 203931 194024 203959
rect 193864 203897 194024 203931
rect 193864 203869 193899 203897
rect 193927 203869 193961 203897
rect 193989 203869 194024 203897
rect 193864 203835 194024 203869
rect 193864 203807 193899 203835
rect 193927 203807 193961 203835
rect 193989 203807 194024 203835
rect 193864 203773 194024 203807
rect 193864 203745 193899 203773
rect 193927 203745 193961 203773
rect 193989 203745 194024 203773
rect 193864 203728 194024 203745
rect 209224 203959 209384 203976
rect 209224 203931 209259 203959
rect 209287 203931 209321 203959
rect 209349 203931 209384 203959
rect 209224 203897 209384 203931
rect 209224 203869 209259 203897
rect 209287 203869 209321 203897
rect 209349 203869 209384 203897
rect 209224 203835 209384 203869
rect 209224 203807 209259 203835
rect 209287 203807 209321 203835
rect 209349 203807 209384 203835
rect 209224 203773 209384 203807
rect 209224 203745 209259 203773
rect 209287 203745 209321 203773
rect 209349 203745 209384 203773
rect 209224 203728 209384 203745
rect 224584 203959 224744 203976
rect 224584 203931 224619 203959
rect 224647 203931 224681 203959
rect 224709 203931 224744 203959
rect 224584 203897 224744 203931
rect 224584 203869 224619 203897
rect 224647 203869 224681 203897
rect 224709 203869 224744 203897
rect 224584 203835 224744 203869
rect 224584 203807 224619 203835
rect 224647 203807 224681 203835
rect 224709 203807 224744 203835
rect 224584 203773 224744 203807
rect 224584 203745 224619 203773
rect 224647 203745 224681 203773
rect 224709 203745 224744 203773
rect 224584 203728 224744 203745
rect 239944 203959 240104 203976
rect 239944 203931 239979 203959
rect 240007 203931 240041 203959
rect 240069 203931 240104 203959
rect 239944 203897 240104 203931
rect 239944 203869 239979 203897
rect 240007 203869 240041 203897
rect 240069 203869 240104 203897
rect 239944 203835 240104 203869
rect 239944 203807 239979 203835
rect 240007 203807 240041 203835
rect 240069 203807 240104 203835
rect 239944 203773 240104 203807
rect 239944 203745 239979 203773
rect 240007 203745 240041 203773
rect 240069 203745 240104 203773
rect 239944 203728 240104 203745
rect 32584 200959 32744 200976
rect 32584 200931 32619 200959
rect 32647 200931 32681 200959
rect 32709 200931 32744 200959
rect 32584 200897 32744 200931
rect 32584 200869 32619 200897
rect 32647 200869 32681 200897
rect 32709 200869 32744 200897
rect 32584 200835 32744 200869
rect 32584 200807 32619 200835
rect 32647 200807 32681 200835
rect 32709 200807 32744 200835
rect 32584 200773 32744 200807
rect 32584 200745 32619 200773
rect 32647 200745 32681 200773
rect 32709 200745 32744 200773
rect 32584 200728 32744 200745
rect 47944 200959 48104 200976
rect 47944 200931 47979 200959
rect 48007 200931 48041 200959
rect 48069 200931 48104 200959
rect 47944 200897 48104 200931
rect 47944 200869 47979 200897
rect 48007 200869 48041 200897
rect 48069 200869 48104 200897
rect 47944 200835 48104 200869
rect 47944 200807 47979 200835
rect 48007 200807 48041 200835
rect 48069 200807 48104 200835
rect 47944 200773 48104 200807
rect 47944 200745 47979 200773
rect 48007 200745 48041 200773
rect 48069 200745 48104 200773
rect 47944 200728 48104 200745
rect 63304 200959 63464 200976
rect 63304 200931 63339 200959
rect 63367 200931 63401 200959
rect 63429 200931 63464 200959
rect 63304 200897 63464 200931
rect 63304 200869 63339 200897
rect 63367 200869 63401 200897
rect 63429 200869 63464 200897
rect 63304 200835 63464 200869
rect 63304 200807 63339 200835
rect 63367 200807 63401 200835
rect 63429 200807 63464 200835
rect 63304 200773 63464 200807
rect 63304 200745 63339 200773
rect 63367 200745 63401 200773
rect 63429 200745 63464 200773
rect 63304 200728 63464 200745
rect 78664 200959 78824 200976
rect 78664 200931 78699 200959
rect 78727 200931 78761 200959
rect 78789 200931 78824 200959
rect 78664 200897 78824 200931
rect 78664 200869 78699 200897
rect 78727 200869 78761 200897
rect 78789 200869 78824 200897
rect 78664 200835 78824 200869
rect 78664 200807 78699 200835
rect 78727 200807 78761 200835
rect 78789 200807 78824 200835
rect 78664 200773 78824 200807
rect 78664 200745 78699 200773
rect 78727 200745 78761 200773
rect 78789 200745 78824 200773
rect 78664 200728 78824 200745
rect 94024 200959 94184 200976
rect 94024 200931 94059 200959
rect 94087 200931 94121 200959
rect 94149 200931 94184 200959
rect 94024 200897 94184 200931
rect 94024 200869 94059 200897
rect 94087 200869 94121 200897
rect 94149 200869 94184 200897
rect 94024 200835 94184 200869
rect 94024 200807 94059 200835
rect 94087 200807 94121 200835
rect 94149 200807 94184 200835
rect 94024 200773 94184 200807
rect 94024 200745 94059 200773
rect 94087 200745 94121 200773
rect 94149 200745 94184 200773
rect 94024 200728 94184 200745
rect 109384 200959 109544 200976
rect 109384 200931 109419 200959
rect 109447 200931 109481 200959
rect 109509 200931 109544 200959
rect 109384 200897 109544 200931
rect 109384 200869 109419 200897
rect 109447 200869 109481 200897
rect 109509 200869 109544 200897
rect 109384 200835 109544 200869
rect 109384 200807 109419 200835
rect 109447 200807 109481 200835
rect 109509 200807 109544 200835
rect 109384 200773 109544 200807
rect 109384 200745 109419 200773
rect 109447 200745 109481 200773
rect 109509 200745 109544 200773
rect 109384 200728 109544 200745
rect 124744 200959 124904 200976
rect 124744 200931 124779 200959
rect 124807 200931 124841 200959
rect 124869 200931 124904 200959
rect 124744 200897 124904 200931
rect 124744 200869 124779 200897
rect 124807 200869 124841 200897
rect 124869 200869 124904 200897
rect 124744 200835 124904 200869
rect 124744 200807 124779 200835
rect 124807 200807 124841 200835
rect 124869 200807 124904 200835
rect 124744 200773 124904 200807
rect 124744 200745 124779 200773
rect 124807 200745 124841 200773
rect 124869 200745 124904 200773
rect 124744 200728 124904 200745
rect 140104 200959 140264 200976
rect 140104 200931 140139 200959
rect 140167 200931 140201 200959
rect 140229 200931 140264 200959
rect 140104 200897 140264 200931
rect 140104 200869 140139 200897
rect 140167 200869 140201 200897
rect 140229 200869 140264 200897
rect 140104 200835 140264 200869
rect 140104 200807 140139 200835
rect 140167 200807 140201 200835
rect 140229 200807 140264 200835
rect 140104 200773 140264 200807
rect 140104 200745 140139 200773
rect 140167 200745 140201 200773
rect 140229 200745 140264 200773
rect 140104 200728 140264 200745
rect 155464 200959 155624 200976
rect 155464 200931 155499 200959
rect 155527 200931 155561 200959
rect 155589 200931 155624 200959
rect 155464 200897 155624 200931
rect 155464 200869 155499 200897
rect 155527 200869 155561 200897
rect 155589 200869 155624 200897
rect 155464 200835 155624 200869
rect 155464 200807 155499 200835
rect 155527 200807 155561 200835
rect 155589 200807 155624 200835
rect 155464 200773 155624 200807
rect 155464 200745 155499 200773
rect 155527 200745 155561 200773
rect 155589 200745 155624 200773
rect 155464 200728 155624 200745
rect 170824 200959 170984 200976
rect 170824 200931 170859 200959
rect 170887 200931 170921 200959
rect 170949 200931 170984 200959
rect 170824 200897 170984 200931
rect 170824 200869 170859 200897
rect 170887 200869 170921 200897
rect 170949 200869 170984 200897
rect 170824 200835 170984 200869
rect 170824 200807 170859 200835
rect 170887 200807 170921 200835
rect 170949 200807 170984 200835
rect 170824 200773 170984 200807
rect 170824 200745 170859 200773
rect 170887 200745 170921 200773
rect 170949 200745 170984 200773
rect 170824 200728 170984 200745
rect 186184 200959 186344 200976
rect 186184 200931 186219 200959
rect 186247 200931 186281 200959
rect 186309 200931 186344 200959
rect 186184 200897 186344 200931
rect 186184 200869 186219 200897
rect 186247 200869 186281 200897
rect 186309 200869 186344 200897
rect 186184 200835 186344 200869
rect 186184 200807 186219 200835
rect 186247 200807 186281 200835
rect 186309 200807 186344 200835
rect 186184 200773 186344 200807
rect 186184 200745 186219 200773
rect 186247 200745 186281 200773
rect 186309 200745 186344 200773
rect 186184 200728 186344 200745
rect 201544 200959 201704 200976
rect 201544 200931 201579 200959
rect 201607 200931 201641 200959
rect 201669 200931 201704 200959
rect 201544 200897 201704 200931
rect 201544 200869 201579 200897
rect 201607 200869 201641 200897
rect 201669 200869 201704 200897
rect 201544 200835 201704 200869
rect 201544 200807 201579 200835
rect 201607 200807 201641 200835
rect 201669 200807 201704 200835
rect 201544 200773 201704 200807
rect 201544 200745 201579 200773
rect 201607 200745 201641 200773
rect 201669 200745 201704 200773
rect 201544 200728 201704 200745
rect 216904 200959 217064 200976
rect 216904 200931 216939 200959
rect 216967 200931 217001 200959
rect 217029 200931 217064 200959
rect 216904 200897 217064 200931
rect 216904 200869 216939 200897
rect 216967 200869 217001 200897
rect 217029 200869 217064 200897
rect 216904 200835 217064 200869
rect 216904 200807 216939 200835
rect 216967 200807 217001 200835
rect 217029 200807 217064 200835
rect 216904 200773 217064 200807
rect 216904 200745 216939 200773
rect 216967 200745 217001 200773
rect 217029 200745 217064 200773
rect 216904 200728 217064 200745
rect 232264 200959 232424 200976
rect 232264 200931 232299 200959
rect 232327 200931 232361 200959
rect 232389 200931 232424 200959
rect 232264 200897 232424 200931
rect 232264 200869 232299 200897
rect 232327 200869 232361 200897
rect 232389 200869 232424 200897
rect 232264 200835 232424 200869
rect 232264 200807 232299 200835
rect 232327 200807 232361 200835
rect 232389 200807 232424 200835
rect 232264 200773 232424 200807
rect 232264 200745 232299 200773
rect 232327 200745 232361 200773
rect 232389 200745 232424 200773
rect 232264 200728 232424 200745
rect 247624 200959 247784 200976
rect 247624 200931 247659 200959
rect 247687 200931 247721 200959
rect 247749 200931 247784 200959
rect 247624 200897 247784 200931
rect 247624 200869 247659 200897
rect 247687 200869 247721 200897
rect 247749 200869 247784 200897
rect 247624 200835 247784 200869
rect 247624 200807 247659 200835
rect 247687 200807 247721 200835
rect 247749 200807 247784 200835
rect 247624 200773 247784 200807
rect 247624 200745 247659 200773
rect 247687 200745 247721 200773
rect 247749 200745 247784 200773
rect 247624 200728 247784 200745
rect 254529 200959 254839 209745
rect 254529 200931 254577 200959
rect 254605 200931 254639 200959
rect 254667 200931 254701 200959
rect 254729 200931 254763 200959
rect 254791 200931 254839 200959
rect 254529 200897 254839 200931
rect 254529 200869 254577 200897
rect 254605 200869 254639 200897
rect 254667 200869 254701 200897
rect 254729 200869 254763 200897
rect 254791 200869 254839 200897
rect 254529 200835 254839 200869
rect 254529 200807 254577 200835
rect 254605 200807 254639 200835
rect 254667 200807 254701 200835
rect 254729 200807 254763 200835
rect 254791 200807 254839 200835
rect 254529 200773 254839 200807
rect 254529 200745 254577 200773
rect 254605 200745 254639 200773
rect 254667 200745 254701 200773
rect 254729 200745 254763 200773
rect 254791 200745 254839 200773
rect 31389 194931 31437 194959
rect 31465 194931 31499 194959
rect 31527 194931 31561 194959
rect 31589 194931 31623 194959
rect 31651 194931 31699 194959
rect 31389 194897 31699 194931
rect 31389 194869 31437 194897
rect 31465 194869 31499 194897
rect 31527 194869 31561 194897
rect 31589 194869 31623 194897
rect 31651 194869 31699 194897
rect 31389 194835 31699 194869
rect 31389 194807 31437 194835
rect 31465 194807 31499 194835
rect 31527 194807 31561 194835
rect 31589 194807 31623 194835
rect 31651 194807 31699 194835
rect 31389 194773 31699 194807
rect 31389 194745 31437 194773
rect 31465 194745 31499 194773
rect 31527 194745 31561 194773
rect 31589 194745 31623 194773
rect 31651 194745 31699 194773
rect 31389 185959 31699 194745
rect 40264 194959 40424 194976
rect 40264 194931 40299 194959
rect 40327 194931 40361 194959
rect 40389 194931 40424 194959
rect 40264 194897 40424 194931
rect 40264 194869 40299 194897
rect 40327 194869 40361 194897
rect 40389 194869 40424 194897
rect 40264 194835 40424 194869
rect 40264 194807 40299 194835
rect 40327 194807 40361 194835
rect 40389 194807 40424 194835
rect 40264 194773 40424 194807
rect 40264 194745 40299 194773
rect 40327 194745 40361 194773
rect 40389 194745 40424 194773
rect 40264 194728 40424 194745
rect 55624 194959 55784 194976
rect 55624 194931 55659 194959
rect 55687 194931 55721 194959
rect 55749 194931 55784 194959
rect 55624 194897 55784 194931
rect 55624 194869 55659 194897
rect 55687 194869 55721 194897
rect 55749 194869 55784 194897
rect 55624 194835 55784 194869
rect 55624 194807 55659 194835
rect 55687 194807 55721 194835
rect 55749 194807 55784 194835
rect 55624 194773 55784 194807
rect 55624 194745 55659 194773
rect 55687 194745 55721 194773
rect 55749 194745 55784 194773
rect 55624 194728 55784 194745
rect 70984 194959 71144 194976
rect 70984 194931 71019 194959
rect 71047 194931 71081 194959
rect 71109 194931 71144 194959
rect 70984 194897 71144 194931
rect 70984 194869 71019 194897
rect 71047 194869 71081 194897
rect 71109 194869 71144 194897
rect 70984 194835 71144 194869
rect 70984 194807 71019 194835
rect 71047 194807 71081 194835
rect 71109 194807 71144 194835
rect 70984 194773 71144 194807
rect 70984 194745 71019 194773
rect 71047 194745 71081 194773
rect 71109 194745 71144 194773
rect 70984 194728 71144 194745
rect 86344 194959 86504 194976
rect 86344 194931 86379 194959
rect 86407 194931 86441 194959
rect 86469 194931 86504 194959
rect 86344 194897 86504 194931
rect 86344 194869 86379 194897
rect 86407 194869 86441 194897
rect 86469 194869 86504 194897
rect 86344 194835 86504 194869
rect 86344 194807 86379 194835
rect 86407 194807 86441 194835
rect 86469 194807 86504 194835
rect 86344 194773 86504 194807
rect 86344 194745 86379 194773
rect 86407 194745 86441 194773
rect 86469 194745 86504 194773
rect 86344 194728 86504 194745
rect 101704 194959 101864 194976
rect 101704 194931 101739 194959
rect 101767 194931 101801 194959
rect 101829 194931 101864 194959
rect 101704 194897 101864 194931
rect 101704 194869 101739 194897
rect 101767 194869 101801 194897
rect 101829 194869 101864 194897
rect 101704 194835 101864 194869
rect 101704 194807 101739 194835
rect 101767 194807 101801 194835
rect 101829 194807 101864 194835
rect 101704 194773 101864 194807
rect 101704 194745 101739 194773
rect 101767 194745 101801 194773
rect 101829 194745 101864 194773
rect 101704 194728 101864 194745
rect 117064 194959 117224 194976
rect 117064 194931 117099 194959
rect 117127 194931 117161 194959
rect 117189 194931 117224 194959
rect 117064 194897 117224 194931
rect 117064 194869 117099 194897
rect 117127 194869 117161 194897
rect 117189 194869 117224 194897
rect 117064 194835 117224 194869
rect 117064 194807 117099 194835
rect 117127 194807 117161 194835
rect 117189 194807 117224 194835
rect 117064 194773 117224 194807
rect 117064 194745 117099 194773
rect 117127 194745 117161 194773
rect 117189 194745 117224 194773
rect 117064 194728 117224 194745
rect 132424 194959 132584 194976
rect 132424 194931 132459 194959
rect 132487 194931 132521 194959
rect 132549 194931 132584 194959
rect 132424 194897 132584 194931
rect 132424 194869 132459 194897
rect 132487 194869 132521 194897
rect 132549 194869 132584 194897
rect 132424 194835 132584 194869
rect 132424 194807 132459 194835
rect 132487 194807 132521 194835
rect 132549 194807 132584 194835
rect 132424 194773 132584 194807
rect 132424 194745 132459 194773
rect 132487 194745 132521 194773
rect 132549 194745 132584 194773
rect 132424 194728 132584 194745
rect 147784 194959 147944 194976
rect 147784 194931 147819 194959
rect 147847 194931 147881 194959
rect 147909 194931 147944 194959
rect 147784 194897 147944 194931
rect 147784 194869 147819 194897
rect 147847 194869 147881 194897
rect 147909 194869 147944 194897
rect 147784 194835 147944 194869
rect 147784 194807 147819 194835
rect 147847 194807 147881 194835
rect 147909 194807 147944 194835
rect 147784 194773 147944 194807
rect 147784 194745 147819 194773
rect 147847 194745 147881 194773
rect 147909 194745 147944 194773
rect 147784 194728 147944 194745
rect 163144 194959 163304 194976
rect 163144 194931 163179 194959
rect 163207 194931 163241 194959
rect 163269 194931 163304 194959
rect 163144 194897 163304 194931
rect 163144 194869 163179 194897
rect 163207 194869 163241 194897
rect 163269 194869 163304 194897
rect 163144 194835 163304 194869
rect 163144 194807 163179 194835
rect 163207 194807 163241 194835
rect 163269 194807 163304 194835
rect 163144 194773 163304 194807
rect 163144 194745 163179 194773
rect 163207 194745 163241 194773
rect 163269 194745 163304 194773
rect 163144 194728 163304 194745
rect 178504 194959 178664 194976
rect 178504 194931 178539 194959
rect 178567 194931 178601 194959
rect 178629 194931 178664 194959
rect 178504 194897 178664 194931
rect 178504 194869 178539 194897
rect 178567 194869 178601 194897
rect 178629 194869 178664 194897
rect 178504 194835 178664 194869
rect 178504 194807 178539 194835
rect 178567 194807 178601 194835
rect 178629 194807 178664 194835
rect 178504 194773 178664 194807
rect 178504 194745 178539 194773
rect 178567 194745 178601 194773
rect 178629 194745 178664 194773
rect 178504 194728 178664 194745
rect 193864 194959 194024 194976
rect 193864 194931 193899 194959
rect 193927 194931 193961 194959
rect 193989 194931 194024 194959
rect 193864 194897 194024 194931
rect 193864 194869 193899 194897
rect 193927 194869 193961 194897
rect 193989 194869 194024 194897
rect 193864 194835 194024 194869
rect 193864 194807 193899 194835
rect 193927 194807 193961 194835
rect 193989 194807 194024 194835
rect 193864 194773 194024 194807
rect 193864 194745 193899 194773
rect 193927 194745 193961 194773
rect 193989 194745 194024 194773
rect 193864 194728 194024 194745
rect 209224 194959 209384 194976
rect 209224 194931 209259 194959
rect 209287 194931 209321 194959
rect 209349 194931 209384 194959
rect 209224 194897 209384 194931
rect 209224 194869 209259 194897
rect 209287 194869 209321 194897
rect 209349 194869 209384 194897
rect 209224 194835 209384 194869
rect 209224 194807 209259 194835
rect 209287 194807 209321 194835
rect 209349 194807 209384 194835
rect 209224 194773 209384 194807
rect 209224 194745 209259 194773
rect 209287 194745 209321 194773
rect 209349 194745 209384 194773
rect 209224 194728 209384 194745
rect 224584 194959 224744 194976
rect 224584 194931 224619 194959
rect 224647 194931 224681 194959
rect 224709 194931 224744 194959
rect 224584 194897 224744 194931
rect 224584 194869 224619 194897
rect 224647 194869 224681 194897
rect 224709 194869 224744 194897
rect 224584 194835 224744 194869
rect 224584 194807 224619 194835
rect 224647 194807 224681 194835
rect 224709 194807 224744 194835
rect 224584 194773 224744 194807
rect 224584 194745 224619 194773
rect 224647 194745 224681 194773
rect 224709 194745 224744 194773
rect 224584 194728 224744 194745
rect 239944 194959 240104 194976
rect 239944 194931 239979 194959
rect 240007 194931 240041 194959
rect 240069 194931 240104 194959
rect 239944 194897 240104 194931
rect 239944 194869 239979 194897
rect 240007 194869 240041 194897
rect 240069 194869 240104 194897
rect 239944 194835 240104 194869
rect 239944 194807 239979 194835
rect 240007 194807 240041 194835
rect 240069 194807 240104 194835
rect 239944 194773 240104 194807
rect 239944 194745 239979 194773
rect 240007 194745 240041 194773
rect 240069 194745 240104 194773
rect 239944 194728 240104 194745
rect 32584 191959 32744 191976
rect 32584 191931 32619 191959
rect 32647 191931 32681 191959
rect 32709 191931 32744 191959
rect 32584 191897 32744 191931
rect 32584 191869 32619 191897
rect 32647 191869 32681 191897
rect 32709 191869 32744 191897
rect 32584 191835 32744 191869
rect 32584 191807 32619 191835
rect 32647 191807 32681 191835
rect 32709 191807 32744 191835
rect 32584 191773 32744 191807
rect 32584 191745 32619 191773
rect 32647 191745 32681 191773
rect 32709 191745 32744 191773
rect 32584 191728 32744 191745
rect 47944 191959 48104 191976
rect 47944 191931 47979 191959
rect 48007 191931 48041 191959
rect 48069 191931 48104 191959
rect 47944 191897 48104 191931
rect 47944 191869 47979 191897
rect 48007 191869 48041 191897
rect 48069 191869 48104 191897
rect 47944 191835 48104 191869
rect 47944 191807 47979 191835
rect 48007 191807 48041 191835
rect 48069 191807 48104 191835
rect 47944 191773 48104 191807
rect 47944 191745 47979 191773
rect 48007 191745 48041 191773
rect 48069 191745 48104 191773
rect 47944 191728 48104 191745
rect 63304 191959 63464 191976
rect 63304 191931 63339 191959
rect 63367 191931 63401 191959
rect 63429 191931 63464 191959
rect 63304 191897 63464 191931
rect 63304 191869 63339 191897
rect 63367 191869 63401 191897
rect 63429 191869 63464 191897
rect 63304 191835 63464 191869
rect 63304 191807 63339 191835
rect 63367 191807 63401 191835
rect 63429 191807 63464 191835
rect 63304 191773 63464 191807
rect 63304 191745 63339 191773
rect 63367 191745 63401 191773
rect 63429 191745 63464 191773
rect 63304 191728 63464 191745
rect 78664 191959 78824 191976
rect 78664 191931 78699 191959
rect 78727 191931 78761 191959
rect 78789 191931 78824 191959
rect 78664 191897 78824 191931
rect 78664 191869 78699 191897
rect 78727 191869 78761 191897
rect 78789 191869 78824 191897
rect 78664 191835 78824 191869
rect 78664 191807 78699 191835
rect 78727 191807 78761 191835
rect 78789 191807 78824 191835
rect 78664 191773 78824 191807
rect 78664 191745 78699 191773
rect 78727 191745 78761 191773
rect 78789 191745 78824 191773
rect 78664 191728 78824 191745
rect 94024 191959 94184 191976
rect 94024 191931 94059 191959
rect 94087 191931 94121 191959
rect 94149 191931 94184 191959
rect 94024 191897 94184 191931
rect 94024 191869 94059 191897
rect 94087 191869 94121 191897
rect 94149 191869 94184 191897
rect 94024 191835 94184 191869
rect 94024 191807 94059 191835
rect 94087 191807 94121 191835
rect 94149 191807 94184 191835
rect 94024 191773 94184 191807
rect 94024 191745 94059 191773
rect 94087 191745 94121 191773
rect 94149 191745 94184 191773
rect 94024 191728 94184 191745
rect 109384 191959 109544 191976
rect 109384 191931 109419 191959
rect 109447 191931 109481 191959
rect 109509 191931 109544 191959
rect 109384 191897 109544 191931
rect 109384 191869 109419 191897
rect 109447 191869 109481 191897
rect 109509 191869 109544 191897
rect 109384 191835 109544 191869
rect 109384 191807 109419 191835
rect 109447 191807 109481 191835
rect 109509 191807 109544 191835
rect 109384 191773 109544 191807
rect 109384 191745 109419 191773
rect 109447 191745 109481 191773
rect 109509 191745 109544 191773
rect 109384 191728 109544 191745
rect 124744 191959 124904 191976
rect 124744 191931 124779 191959
rect 124807 191931 124841 191959
rect 124869 191931 124904 191959
rect 124744 191897 124904 191931
rect 124744 191869 124779 191897
rect 124807 191869 124841 191897
rect 124869 191869 124904 191897
rect 124744 191835 124904 191869
rect 124744 191807 124779 191835
rect 124807 191807 124841 191835
rect 124869 191807 124904 191835
rect 124744 191773 124904 191807
rect 124744 191745 124779 191773
rect 124807 191745 124841 191773
rect 124869 191745 124904 191773
rect 124744 191728 124904 191745
rect 140104 191959 140264 191976
rect 140104 191931 140139 191959
rect 140167 191931 140201 191959
rect 140229 191931 140264 191959
rect 140104 191897 140264 191931
rect 140104 191869 140139 191897
rect 140167 191869 140201 191897
rect 140229 191869 140264 191897
rect 140104 191835 140264 191869
rect 140104 191807 140139 191835
rect 140167 191807 140201 191835
rect 140229 191807 140264 191835
rect 140104 191773 140264 191807
rect 140104 191745 140139 191773
rect 140167 191745 140201 191773
rect 140229 191745 140264 191773
rect 140104 191728 140264 191745
rect 155464 191959 155624 191976
rect 155464 191931 155499 191959
rect 155527 191931 155561 191959
rect 155589 191931 155624 191959
rect 155464 191897 155624 191931
rect 155464 191869 155499 191897
rect 155527 191869 155561 191897
rect 155589 191869 155624 191897
rect 155464 191835 155624 191869
rect 155464 191807 155499 191835
rect 155527 191807 155561 191835
rect 155589 191807 155624 191835
rect 155464 191773 155624 191807
rect 155464 191745 155499 191773
rect 155527 191745 155561 191773
rect 155589 191745 155624 191773
rect 155464 191728 155624 191745
rect 170824 191959 170984 191976
rect 170824 191931 170859 191959
rect 170887 191931 170921 191959
rect 170949 191931 170984 191959
rect 170824 191897 170984 191931
rect 170824 191869 170859 191897
rect 170887 191869 170921 191897
rect 170949 191869 170984 191897
rect 170824 191835 170984 191869
rect 170824 191807 170859 191835
rect 170887 191807 170921 191835
rect 170949 191807 170984 191835
rect 170824 191773 170984 191807
rect 170824 191745 170859 191773
rect 170887 191745 170921 191773
rect 170949 191745 170984 191773
rect 170824 191728 170984 191745
rect 186184 191959 186344 191976
rect 186184 191931 186219 191959
rect 186247 191931 186281 191959
rect 186309 191931 186344 191959
rect 186184 191897 186344 191931
rect 186184 191869 186219 191897
rect 186247 191869 186281 191897
rect 186309 191869 186344 191897
rect 186184 191835 186344 191869
rect 186184 191807 186219 191835
rect 186247 191807 186281 191835
rect 186309 191807 186344 191835
rect 186184 191773 186344 191807
rect 186184 191745 186219 191773
rect 186247 191745 186281 191773
rect 186309 191745 186344 191773
rect 186184 191728 186344 191745
rect 201544 191959 201704 191976
rect 201544 191931 201579 191959
rect 201607 191931 201641 191959
rect 201669 191931 201704 191959
rect 201544 191897 201704 191931
rect 201544 191869 201579 191897
rect 201607 191869 201641 191897
rect 201669 191869 201704 191897
rect 201544 191835 201704 191869
rect 201544 191807 201579 191835
rect 201607 191807 201641 191835
rect 201669 191807 201704 191835
rect 201544 191773 201704 191807
rect 201544 191745 201579 191773
rect 201607 191745 201641 191773
rect 201669 191745 201704 191773
rect 201544 191728 201704 191745
rect 216904 191959 217064 191976
rect 216904 191931 216939 191959
rect 216967 191931 217001 191959
rect 217029 191931 217064 191959
rect 216904 191897 217064 191931
rect 216904 191869 216939 191897
rect 216967 191869 217001 191897
rect 217029 191869 217064 191897
rect 216904 191835 217064 191869
rect 216904 191807 216939 191835
rect 216967 191807 217001 191835
rect 217029 191807 217064 191835
rect 216904 191773 217064 191807
rect 216904 191745 216939 191773
rect 216967 191745 217001 191773
rect 217029 191745 217064 191773
rect 216904 191728 217064 191745
rect 232264 191959 232424 191976
rect 232264 191931 232299 191959
rect 232327 191931 232361 191959
rect 232389 191931 232424 191959
rect 232264 191897 232424 191931
rect 232264 191869 232299 191897
rect 232327 191869 232361 191897
rect 232389 191869 232424 191897
rect 232264 191835 232424 191869
rect 232264 191807 232299 191835
rect 232327 191807 232361 191835
rect 232389 191807 232424 191835
rect 232264 191773 232424 191807
rect 232264 191745 232299 191773
rect 232327 191745 232361 191773
rect 232389 191745 232424 191773
rect 232264 191728 232424 191745
rect 247624 191959 247784 191976
rect 247624 191931 247659 191959
rect 247687 191931 247721 191959
rect 247749 191931 247784 191959
rect 247624 191897 247784 191931
rect 247624 191869 247659 191897
rect 247687 191869 247721 191897
rect 247749 191869 247784 191897
rect 247624 191835 247784 191869
rect 247624 191807 247659 191835
rect 247687 191807 247721 191835
rect 247749 191807 247784 191835
rect 247624 191773 247784 191807
rect 247624 191745 247659 191773
rect 247687 191745 247721 191773
rect 247749 191745 247784 191773
rect 247624 191728 247784 191745
rect 254529 191959 254839 200745
rect 254529 191931 254577 191959
rect 254605 191931 254639 191959
rect 254667 191931 254701 191959
rect 254729 191931 254763 191959
rect 254791 191931 254839 191959
rect 254529 191897 254839 191931
rect 254529 191869 254577 191897
rect 254605 191869 254639 191897
rect 254667 191869 254701 191897
rect 254729 191869 254763 191897
rect 254791 191869 254839 191897
rect 254529 191835 254839 191869
rect 254529 191807 254577 191835
rect 254605 191807 254639 191835
rect 254667 191807 254701 191835
rect 254729 191807 254763 191835
rect 254791 191807 254839 191835
rect 254529 191773 254839 191807
rect 254529 191745 254577 191773
rect 254605 191745 254639 191773
rect 254667 191745 254701 191773
rect 254729 191745 254763 191773
rect 254791 191745 254839 191773
rect 31389 185931 31437 185959
rect 31465 185931 31499 185959
rect 31527 185931 31561 185959
rect 31589 185931 31623 185959
rect 31651 185931 31699 185959
rect 31389 185897 31699 185931
rect 31389 185869 31437 185897
rect 31465 185869 31499 185897
rect 31527 185869 31561 185897
rect 31589 185869 31623 185897
rect 31651 185869 31699 185897
rect 31389 185835 31699 185869
rect 31389 185807 31437 185835
rect 31465 185807 31499 185835
rect 31527 185807 31561 185835
rect 31589 185807 31623 185835
rect 31651 185807 31699 185835
rect 31389 185773 31699 185807
rect 31389 185745 31437 185773
rect 31465 185745 31499 185773
rect 31527 185745 31561 185773
rect 31589 185745 31623 185773
rect 31651 185745 31699 185773
rect 31389 176959 31699 185745
rect 40264 185959 40424 185976
rect 40264 185931 40299 185959
rect 40327 185931 40361 185959
rect 40389 185931 40424 185959
rect 40264 185897 40424 185931
rect 40264 185869 40299 185897
rect 40327 185869 40361 185897
rect 40389 185869 40424 185897
rect 40264 185835 40424 185869
rect 40264 185807 40299 185835
rect 40327 185807 40361 185835
rect 40389 185807 40424 185835
rect 40264 185773 40424 185807
rect 40264 185745 40299 185773
rect 40327 185745 40361 185773
rect 40389 185745 40424 185773
rect 40264 185728 40424 185745
rect 55624 185959 55784 185976
rect 55624 185931 55659 185959
rect 55687 185931 55721 185959
rect 55749 185931 55784 185959
rect 55624 185897 55784 185931
rect 55624 185869 55659 185897
rect 55687 185869 55721 185897
rect 55749 185869 55784 185897
rect 55624 185835 55784 185869
rect 55624 185807 55659 185835
rect 55687 185807 55721 185835
rect 55749 185807 55784 185835
rect 55624 185773 55784 185807
rect 55624 185745 55659 185773
rect 55687 185745 55721 185773
rect 55749 185745 55784 185773
rect 55624 185728 55784 185745
rect 70984 185959 71144 185976
rect 70984 185931 71019 185959
rect 71047 185931 71081 185959
rect 71109 185931 71144 185959
rect 70984 185897 71144 185931
rect 70984 185869 71019 185897
rect 71047 185869 71081 185897
rect 71109 185869 71144 185897
rect 70984 185835 71144 185869
rect 70984 185807 71019 185835
rect 71047 185807 71081 185835
rect 71109 185807 71144 185835
rect 70984 185773 71144 185807
rect 70984 185745 71019 185773
rect 71047 185745 71081 185773
rect 71109 185745 71144 185773
rect 70984 185728 71144 185745
rect 86344 185959 86504 185976
rect 86344 185931 86379 185959
rect 86407 185931 86441 185959
rect 86469 185931 86504 185959
rect 86344 185897 86504 185931
rect 86344 185869 86379 185897
rect 86407 185869 86441 185897
rect 86469 185869 86504 185897
rect 86344 185835 86504 185869
rect 86344 185807 86379 185835
rect 86407 185807 86441 185835
rect 86469 185807 86504 185835
rect 86344 185773 86504 185807
rect 86344 185745 86379 185773
rect 86407 185745 86441 185773
rect 86469 185745 86504 185773
rect 86344 185728 86504 185745
rect 101704 185959 101864 185976
rect 101704 185931 101739 185959
rect 101767 185931 101801 185959
rect 101829 185931 101864 185959
rect 101704 185897 101864 185931
rect 101704 185869 101739 185897
rect 101767 185869 101801 185897
rect 101829 185869 101864 185897
rect 101704 185835 101864 185869
rect 101704 185807 101739 185835
rect 101767 185807 101801 185835
rect 101829 185807 101864 185835
rect 101704 185773 101864 185807
rect 101704 185745 101739 185773
rect 101767 185745 101801 185773
rect 101829 185745 101864 185773
rect 101704 185728 101864 185745
rect 117064 185959 117224 185976
rect 117064 185931 117099 185959
rect 117127 185931 117161 185959
rect 117189 185931 117224 185959
rect 117064 185897 117224 185931
rect 117064 185869 117099 185897
rect 117127 185869 117161 185897
rect 117189 185869 117224 185897
rect 117064 185835 117224 185869
rect 117064 185807 117099 185835
rect 117127 185807 117161 185835
rect 117189 185807 117224 185835
rect 117064 185773 117224 185807
rect 117064 185745 117099 185773
rect 117127 185745 117161 185773
rect 117189 185745 117224 185773
rect 117064 185728 117224 185745
rect 132424 185959 132584 185976
rect 132424 185931 132459 185959
rect 132487 185931 132521 185959
rect 132549 185931 132584 185959
rect 132424 185897 132584 185931
rect 132424 185869 132459 185897
rect 132487 185869 132521 185897
rect 132549 185869 132584 185897
rect 132424 185835 132584 185869
rect 132424 185807 132459 185835
rect 132487 185807 132521 185835
rect 132549 185807 132584 185835
rect 132424 185773 132584 185807
rect 132424 185745 132459 185773
rect 132487 185745 132521 185773
rect 132549 185745 132584 185773
rect 132424 185728 132584 185745
rect 147784 185959 147944 185976
rect 147784 185931 147819 185959
rect 147847 185931 147881 185959
rect 147909 185931 147944 185959
rect 147784 185897 147944 185931
rect 147784 185869 147819 185897
rect 147847 185869 147881 185897
rect 147909 185869 147944 185897
rect 147784 185835 147944 185869
rect 147784 185807 147819 185835
rect 147847 185807 147881 185835
rect 147909 185807 147944 185835
rect 147784 185773 147944 185807
rect 147784 185745 147819 185773
rect 147847 185745 147881 185773
rect 147909 185745 147944 185773
rect 147784 185728 147944 185745
rect 163144 185959 163304 185976
rect 163144 185931 163179 185959
rect 163207 185931 163241 185959
rect 163269 185931 163304 185959
rect 163144 185897 163304 185931
rect 163144 185869 163179 185897
rect 163207 185869 163241 185897
rect 163269 185869 163304 185897
rect 163144 185835 163304 185869
rect 163144 185807 163179 185835
rect 163207 185807 163241 185835
rect 163269 185807 163304 185835
rect 163144 185773 163304 185807
rect 163144 185745 163179 185773
rect 163207 185745 163241 185773
rect 163269 185745 163304 185773
rect 163144 185728 163304 185745
rect 178504 185959 178664 185976
rect 178504 185931 178539 185959
rect 178567 185931 178601 185959
rect 178629 185931 178664 185959
rect 178504 185897 178664 185931
rect 178504 185869 178539 185897
rect 178567 185869 178601 185897
rect 178629 185869 178664 185897
rect 178504 185835 178664 185869
rect 178504 185807 178539 185835
rect 178567 185807 178601 185835
rect 178629 185807 178664 185835
rect 178504 185773 178664 185807
rect 178504 185745 178539 185773
rect 178567 185745 178601 185773
rect 178629 185745 178664 185773
rect 178504 185728 178664 185745
rect 193864 185959 194024 185976
rect 193864 185931 193899 185959
rect 193927 185931 193961 185959
rect 193989 185931 194024 185959
rect 193864 185897 194024 185931
rect 193864 185869 193899 185897
rect 193927 185869 193961 185897
rect 193989 185869 194024 185897
rect 193864 185835 194024 185869
rect 193864 185807 193899 185835
rect 193927 185807 193961 185835
rect 193989 185807 194024 185835
rect 193864 185773 194024 185807
rect 193864 185745 193899 185773
rect 193927 185745 193961 185773
rect 193989 185745 194024 185773
rect 193864 185728 194024 185745
rect 209224 185959 209384 185976
rect 209224 185931 209259 185959
rect 209287 185931 209321 185959
rect 209349 185931 209384 185959
rect 209224 185897 209384 185931
rect 209224 185869 209259 185897
rect 209287 185869 209321 185897
rect 209349 185869 209384 185897
rect 209224 185835 209384 185869
rect 209224 185807 209259 185835
rect 209287 185807 209321 185835
rect 209349 185807 209384 185835
rect 209224 185773 209384 185807
rect 209224 185745 209259 185773
rect 209287 185745 209321 185773
rect 209349 185745 209384 185773
rect 209224 185728 209384 185745
rect 224584 185959 224744 185976
rect 224584 185931 224619 185959
rect 224647 185931 224681 185959
rect 224709 185931 224744 185959
rect 224584 185897 224744 185931
rect 224584 185869 224619 185897
rect 224647 185869 224681 185897
rect 224709 185869 224744 185897
rect 224584 185835 224744 185869
rect 224584 185807 224619 185835
rect 224647 185807 224681 185835
rect 224709 185807 224744 185835
rect 224584 185773 224744 185807
rect 224584 185745 224619 185773
rect 224647 185745 224681 185773
rect 224709 185745 224744 185773
rect 224584 185728 224744 185745
rect 239944 185959 240104 185976
rect 239944 185931 239979 185959
rect 240007 185931 240041 185959
rect 240069 185931 240104 185959
rect 239944 185897 240104 185931
rect 239944 185869 239979 185897
rect 240007 185869 240041 185897
rect 240069 185869 240104 185897
rect 239944 185835 240104 185869
rect 239944 185807 239979 185835
rect 240007 185807 240041 185835
rect 240069 185807 240104 185835
rect 239944 185773 240104 185807
rect 239944 185745 239979 185773
rect 240007 185745 240041 185773
rect 240069 185745 240104 185773
rect 239944 185728 240104 185745
rect 32584 182959 32744 182976
rect 32584 182931 32619 182959
rect 32647 182931 32681 182959
rect 32709 182931 32744 182959
rect 32584 182897 32744 182931
rect 32584 182869 32619 182897
rect 32647 182869 32681 182897
rect 32709 182869 32744 182897
rect 32584 182835 32744 182869
rect 32584 182807 32619 182835
rect 32647 182807 32681 182835
rect 32709 182807 32744 182835
rect 32584 182773 32744 182807
rect 32584 182745 32619 182773
rect 32647 182745 32681 182773
rect 32709 182745 32744 182773
rect 32584 182728 32744 182745
rect 47944 182959 48104 182976
rect 47944 182931 47979 182959
rect 48007 182931 48041 182959
rect 48069 182931 48104 182959
rect 47944 182897 48104 182931
rect 47944 182869 47979 182897
rect 48007 182869 48041 182897
rect 48069 182869 48104 182897
rect 47944 182835 48104 182869
rect 47944 182807 47979 182835
rect 48007 182807 48041 182835
rect 48069 182807 48104 182835
rect 47944 182773 48104 182807
rect 47944 182745 47979 182773
rect 48007 182745 48041 182773
rect 48069 182745 48104 182773
rect 47944 182728 48104 182745
rect 63304 182959 63464 182976
rect 63304 182931 63339 182959
rect 63367 182931 63401 182959
rect 63429 182931 63464 182959
rect 63304 182897 63464 182931
rect 63304 182869 63339 182897
rect 63367 182869 63401 182897
rect 63429 182869 63464 182897
rect 63304 182835 63464 182869
rect 63304 182807 63339 182835
rect 63367 182807 63401 182835
rect 63429 182807 63464 182835
rect 63304 182773 63464 182807
rect 63304 182745 63339 182773
rect 63367 182745 63401 182773
rect 63429 182745 63464 182773
rect 63304 182728 63464 182745
rect 78664 182959 78824 182976
rect 78664 182931 78699 182959
rect 78727 182931 78761 182959
rect 78789 182931 78824 182959
rect 78664 182897 78824 182931
rect 78664 182869 78699 182897
rect 78727 182869 78761 182897
rect 78789 182869 78824 182897
rect 78664 182835 78824 182869
rect 78664 182807 78699 182835
rect 78727 182807 78761 182835
rect 78789 182807 78824 182835
rect 78664 182773 78824 182807
rect 78664 182745 78699 182773
rect 78727 182745 78761 182773
rect 78789 182745 78824 182773
rect 78664 182728 78824 182745
rect 94024 182959 94184 182976
rect 94024 182931 94059 182959
rect 94087 182931 94121 182959
rect 94149 182931 94184 182959
rect 94024 182897 94184 182931
rect 94024 182869 94059 182897
rect 94087 182869 94121 182897
rect 94149 182869 94184 182897
rect 94024 182835 94184 182869
rect 94024 182807 94059 182835
rect 94087 182807 94121 182835
rect 94149 182807 94184 182835
rect 94024 182773 94184 182807
rect 94024 182745 94059 182773
rect 94087 182745 94121 182773
rect 94149 182745 94184 182773
rect 94024 182728 94184 182745
rect 109384 182959 109544 182976
rect 109384 182931 109419 182959
rect 109447 182931 109481 182959
rect 109509 182931 109544 182959
rect 109384 182897 109544 182931
rect 109384 182869 109419 182897
rect 109447 182869 109481 182897
rect 109509 182869 109544 182897
rect 109384 182835 109544 182869
rect 109384 182807 109419 182835
rect 109447 182807 109481 182835
rect 109509 182807 109544 182835
rect 109384 182773 109544 182807
rect 109384 182745 109419 182773
rect 109447 182745 109481 182773
rect 109509 182745 109544 182773
rect 109384 182728 109544 182745
rect 124744 182959 124904 182976
rect 124744 182931 124779 182959
rect 124807 182931 124841 182959
rect 124869 182931 124904 182959
rect 124744 182897 124904 182931
rect 124744 182869 124779 182897
rect 124807 182869 124841 182897
rect 124869 182869 124904 182897
rect 124744 182835 124904 182869
rect 124744 182807 124779 182835
rect 124807 182807 124841 182835
rect 124869 182807 124904 182835
rect 124744 182773 124904 182807
rect 124744 182745 124779 182773
rect 124807 182745 124841 182773
rect 124869 182745 124904 182773
rect 124744 182728 124904 182745
rect 140104 182959 140264 182976
rect 140104 182931 140139 182959
rect 140167 182931 140201 182959
rect 140229 182931 140264 182959
rect 140104 182897 140264 182931
rect 140104 182869 140139 182897
rect 140167 182869 140201 182897
rect 140229 182869 140264 182897
rect 140104 182835 140264 182869
rect 140104 182807 140139 182835
rect 140167 182807 140201 182835
rect 140229 182807 140264 182835
rect 140104 182773 140264 182807
rect 140104 182745 140139 182773
rect 140167 182745 140201 182773
rect 140229 182745 140264 182773
rect 140104 182728 140264 182745
rect 155464 182959 155624 182976
rect 155464 182931 155499 182959
rect 155527 182931 155561 182959
rect 155589 182931 155624 182959
rect 155464 182897 155624 182931
rect 155464 182869 155499 182897
rect 155527 182869 155561 182897
rect 155589 182869 155624 182897
rect 155464 182835 155624 182869
rect 155464 182807 155499 182835
rect 155527 182807 155561 182835
rect 155589 182807 155624 182835
rect 155464 182773 155624 182807
rect 155464 182745 155499 182773
rect 155527 182745 155561 182773
rect 155589 182745 155624 182773
rect 155464 182728 155624 182745
rect 170824 182959 170984 182976
rect 170824 182931 170859 182959
rect 170887 182931 170921 182959
rect 170949 182931 170984 182959
rect 170824 182897 170984 182931
rect 170824 182869 170859 182897
rect 170887 182869 170921 182897
rect 170949 182869 170984 182897
rect 170824 182835 170984 182869
rect 170824 182807 170859 182835
rect 170887 182807 170921 182835
rect 170949 182807 170984 182835
rect 170824 182773 170984 182807
rect 170824 182745 170859 182773
rect 170887 182745 170921 182773
rect 170949 182745 170984 182773
rect 170824 182728 170984 182745
rect 186184 182959 186344 182976
rect 186184 182931 186219 182959
rect 186247 182931 186281 182959
rect 186309 182931 186344 182959
rect 186184 182897 186344 182931
rect 186184 182869 186219 182897
rect 186247 182869 186281 182897
rect 186309 182869 186344 182897
rect 186184 182835 186344 182869
rect 186184 182807 186219 182835
rect 186247 182807 186281 182835
rect 186309 182807 186344 182835
rect 186184 182773 186344 182807
rect 186184 182745 186219 182773
rect 186247 182745 186281 182773
rect 186309 182745 186344 182773
rect 186184 182728 186344 182745
rect 201544 182959 201704 182976
rect 201544 182931 201579 182959
rect 201607 182931 201641 182959
rect 201669 182931 201704 182959
rect 201544 182897 201704 182931
rect 201544 182869 201579 182897
rect 201607 182869 201641 182897
rect 201669 182869 201704 182897
rect 201544 182835 201704 182869
rect 201544 182807 201579 182835
rect 201607 182807 201641 182835
rect 201669 182807 201704 182835
rect 201544 182773 201704 182807
rect 201544 182745 201579 182773
rect 201607 182745 201641 182773
rect 201669 182745 201704 182773
rect 201544 182728 201704 182745
rect 216904 182959 217064 182976
rect 216904 182931 216939 182959
rect 216967 182931 217001 182959
rect 217029 182931 217064 182959
rect 216904 182897 217064 182931
rect 216904 182869 216939 182897
rect 216967 182869 217001 182897
rect 217029 182869 217064 182897
rect 216904 182835 217064 182869
rect 216904 182807 216939 182835
rect 216967 182807 217001 182835
rect 217029 182807 217064 182835
rect 216904 182773 217064 182807
rect 216904 182745 216939 182773
rect 216967 182745 217001 182773
rect 217029 182745 217064 182773
rect 216904 182728 217064 182745
rect 232264 182959 232424 182976
rect 232264 182931 232299 182959
rect 232327 182931 232361 182959
rect 232389 182931 232424 182959
rect 232264 182897 232424 182931
rect 232264 182869 232299 182897
rect 232327 182869 232361 182897
rect 232389 182869 232424 182897
rect 232264 182835 232424 182869
rect 232264 182807 232299 182835
rect 232327 182807 232361 182835
rect 232389 182807 232424 182835
rect 232264 182773 232424 182807
rect 232264 182745 232299 182773
rect 232327 182745 232361 182773
rect 232389 182745 232424 182773
rect 232264 182728 232424 182745
rect 247624 182959 247784 182976
rect 247624 182931 247659 182959
rect 247687 182931 247721 182959
rect 247749 182931 247784 182959
rect 247624 182897 247784 182931
rect 247624 182869 247659 182897
rect 247687 182869 247721 182897
rect 247749 182869 247784 182897
rect 247624 182835 247784 182869
rect 247624 182807 247659 182835
rect 247687 182807 247721 182835
rect 247749 182807 247784 182835
rect 247624 182773 247784 182807
rect 247624 182745 247659 182773
rect 247687 182745 247721 182773
rect 247749 182745 247784 182773
rect 247624 182728 247784 182745
rect 254529 182959 254839 191745
rect 254529 182931 254577 182959
rect 254605 182931 254639 182959
rect 254667 182931 254701 182959
rect 254729 182931 254763 182959
rect 254791 182931 254839 182959
rect 254529 182897 254839 182931
rect 254529 182869 254577 182897
rect 254605 182869 254639 182897
rect 254667 182869 254701 182897
rect 254729 182869 254763 182897
rect 254791 182869 254839 182897
rect 254529 182835 254839 182869
rect 254529 182807 254577 182835
rect 254605 182807 254639 182835
rect 254667 182807 254701 182835
rect 254729 182807 254763 182835
rect 254791 182807 254839 182835
rect 254529 182773 254839 182807
rect 254529 182745 254577 182773
rect 254605 182745 254639 182773
rect 254667 182745 254701 182773
rect 254729 182745 254763 182773
rect 254791 182745 254839 182773
rect 31389 176931 31437 176959
rect 31465 176931 31499 176959
rect 31527 176931 31561 176959
rect 31589 176931 31623 176959
rect 31651 176931 31699 176959
rect 31389 176897 31699 176931
rect 31389 176869 31437 176897
rect 31465 176869 31499 176897
rect 31527 176869 31561 176897
rect 31589 176869 31623 176897
rect 31651 176869 31699 176897
rect 31389 176835 31699 176869
rect 31389 176807 31437 176835
rect 31465 176807 31499 176835
rect 31527 176807 31561 176835
rect 31589 176807 31623 176835
rect 31651 176807 31699 176835
rect 31389 176773 31699 176807
rect 31389 176745 31437 176773
rect 31465 176745 31499 176773
rect 31527 176745 31561 176773
rect 31589 176745 31623 176773
rect 31651 176745 31699 176773
rect 31389 167959 31699 176745
rect 40264 176959 40424 176976
rect 40264 176931 40299 176959
rect 40327 176931 40361 176959
rect 40389 176931 40424 176959
rect 40264 176897 40424 176931
rect 40264 176869 40299 176897
rect 40327 176869 40361 176897
rect 40389 176869 40424 176897
rect 40264 176835 40424 176869
rect 40264 176807 40299 176835
rect 40327 176807 40361 176835
rect 40389 176807 40424 176835
rect 40264 176773 40424 176807
rect 40264 176745 40299 176773
rect 40327 176745 40361 176773
rect 40389 176745 40424 176773
rect 40264 176728 40424 176745
rect 55624 176959 55784 176976
rect 55624 176931 55659 176959
rect 55687 176931 55721 176959
rect 55749 176931 55784 176959
rect 55624 176897 55784 176931
rect 55624 176869 55659 176897
rect 55687 176869 55721 176897
rect 55749 176869 55784 176897
rect 55624 176835 55784 176869
rect 55624 176807 55659 176835
rect 55687 176807 55721 176835
rect 55749 176807 55784 176835
rect 55624 176773 55784 176807
rect 55624 176745 55659 176773
rect 55687 176745 55721 176773
rect 55749 176745 55784 176773
rect 55624 176728 55784 176745
rect 70984 176959 71144 176976
rect 70984 176931 71019 176959
rect 71047 176931 71081 176959
rect 71109 176931 71144 176959
rect 70984 176897 71144 176931
rect 70984 176869 71019 176897
rect 71047 176869 71081 176897
rect 71109 176869 71144 176897
rect 70984 176835 71144 176869
rect 70984 176807 71019 176835
rect 71047 176807 71081 176835
rect 71109 176807 71144 176835
rect 70984 176773 71144 176807
rect 70984 176745 71019 176773
rect 71047 176745 71081 176773
rect 71109 176745 71144 176773
rect 70984 176728 71144 176745
rect 86344 176959 86504 176976
rect 86344 176931 86379 176959
rect 86407 176931 86441 176959
rect 86469 176931 86504 176959
rect 86344 176897 86504 176931
rect 86344 176869 86379 176897
rect 86407 176869 86441 176897
rect 86469 176869 86504 176897
rect 86344 176835 86504 176869
rect 86344 176807 86379 176835
rect 86407 176807 86441 176835
rect 86469 176807 86504 176835
rect 86344 176773 86504 176807
rect 86344 176745 86379 176773
rect 86407 176745 86441 176773
rect 86469 176745 86504 176773
rect 86344 176728 86504 176745
rect 101704 176959 101864 176976
rect 101704 176931 101739 176959
rect 101767 176931 101801 176959
rect 101829 176931 101864 176959
rect 101704 176897 101864 176931
rect 101704 176869 101739 176897
rect 101767 176869 101801 176897
rect 101829 176869 101864 176897
rect 101704 176835 101864 176869
rect 101704 176807 101739 176835
rect 101767 176807 101801 176835
rect 101829 176807 101864 176835
rect 101704 176773 101864 176807
rect 101704 176745 101739 176773
rect 101767 176745 101801 176773
rect 101829 176745 101864 176773
rect 101704 176728 101864 176745
rect 117064 176959 117224 176976
rect 117064 176931 117099 176959
rect 117127 176931 117161 176959
rect 117189 176931 117224 176959
rect 117064 176897 117224 176931
rect 117064 176869 117099 176897
rect 117127 176869 117161 176897
rect 117189 176869 117224 176897
rect 117064 176835 117224 176869
rect 117064 176807 117099 176835
rect 117127 176807 117161 176835
rect 117189 176807 117224 176835
rect 117064 176773 117224 176807
rect 117064 176745 117099 176773
rect 117127 176745 117161 176773
rect 117189 176745 117224 176773
rect 117064 176728 117224 176745
rect 132424 176959 132584 176976
rect 132424 176931 132459 176959
rect 132487 176931 132521 176959
rect 132549 176931 132584 176959
rect 132424 176897 132584 176931
rect 132424 176869 132459 176897
rect 132487 176869 132521 176897
rect 132549 176869 132584 176897
rect 132424 176835 132584 176869
rect 132424 176807 132459 176835
rect 132487 176807 132521 176835
rect 132549 176807 132584 176835
rect 132424 176773 132584 176807
rect 132424 176745 132459 176773
rect 132487 176745 132521 176773
rect 132549 176745 132584 176773
rect 132424 176728 132584 176745
rect 147784 176959 147944 176976
rect 147784 176931 147819 176959
rect 147847 176931 147881 176959
rect 147909 176931 147944 176959
rect 147784 176897 147944 176931
rect 147784 176869 147819 176897
rect 147847 176869 147881 176897
rect 147909 176869 147944 176897
rect 147784 176835 147944 176869
rect 147784 176807 147819 176835
rect 147847 176807 147881 176835
rect 147909 176807 147944 176835
rect 147784 176773 147944 176807
rect 147784 176745 147819 176773
rect 147847 176745 147881 176773
rect 147909 176745 147944 176773
rect 147784 176728 147944 176745
rect 163144 176959 163304 176976
rect 163144 176931 163179 176959
rect 163207 176931 163241 176959
rect 163269 176931 163304 176959
rect 163144 176897 163304 176931
rect 163144 176869 163179 176897
rect 163207 176869 163241 176897
rect 163269 176869 163304 176897
rect 163144 176835 163304 176869
rect 163144 176807 163179 176835
rect 163207 176807 163241 176835
rect 163269 176807 163304 176835
rect 163144 176773 163304 176807
rect 163144 176745 163179 176773
rect 163207 176745 163241 176773
rect 163269 176745 163304 176773
rect 163144 176728 163304 176745
rect 178504 176959 178664 176976
rect 178504 176931 178539 176959
rect 178567 176931 178601 176959
rect 178629 176931 178664 176959
rect 178504 176897 178664 176931
rect 178504 176869 178539 176897
rect 178567 176869 178601 176897
rect 178629 176869 178664 176897
rect 178504 176835 178664 176869
rect 178504 176807 178539 176835
rect 178567 176807 178601 176835
rect 178629 176807 178664 176835
rect 178504 176773 178664 176807
rect 178504 176745 178539 176773
rect 178567 176745 178601 176773
rect 178629 176745 178664 176773
rect 178504 176728 178664 176745
rect 193864 176959 194024 176976
rect 193864 176931 193899 176959
rect 193927 176931 193961 176959
rect 193989 176931 194024 176959
rect 193864 176897 194024 176931
rect 193864 176869 193899 176897
rect 193927 176869 193961 176897
rect 193989 176869 194024 176897
rect 193864 176835 194024 176869
rect 193864 176807 193899 176835
rect 193927 176807 193961 176835
rect 193989 176807 194024 176835
rect 193864 176773 194024 176807
rect 193864 176745 193899 176773
rect 193927 176745 193961 176773
rect 193989 176745 194024 176773
rect 193864 176728 194024 176745
rect 209224 176959 209384 176976
rect 209224 176931 209259 176959
rect 209287 176931 209321 176959
rect 209349 176931 209384 176959
rect 209224 176897 209384 176931
rect 209224 176869 209259 176897
rect 209287 176869 209321 176897
rect 209349 176869 209384 176897
rect 209224 176835 209384 176869
rect 209224 176807 209259 176835
rect 209287 176807 209321 176835
rect 209349 176807 209384 176835
rect 209224 176773 209384 176807
rect 209224 176745 209259 176773
rect 209287 176745 209321 176773
rect 209349 176745 209384 176773
rect 209224 176728 209384 176745
rect 224584 176959 224744 176976
rect 224584 176931 224619 176959
rect 224647 176931 224681 176959
rect 224709 176931 224744 176959
rect 224584 176897 224744 176931
rect 224584 176869 224619 176897
rect 224647 176869 224681 176897
rect 224709 176869 224744 176897
rect 224584 176835 224744 176869
rect 224584 176807 224619 176835
rect 224647 176807 224681 176835
rect 224709 176807 224744 176835
rect 224584 176773 224744 176807
rect 224584 176745 224619 176773
rect 224647 176745 224681 176773
rect 224709 176745 224744 176773
rect 224584 176728 224744 176745
rect 239944 176959 240104 176976
rect 239944 176931 239979 176959
rect 240007 176931 240041 176959
rect 240069 176931 240104 176959
rect 239944 176897 240104 176931
rect 239944 176869 239979 176897
rect 240007 176869 240041 176897
rect 240069 176869 240104 176897
rect 239944 176835 240104 176869
rect 239944 176807 239979 176835
rect 240007 176807 240041 176835
rect 240069 176807 240104 176835
rect 239944 176773 240104 176807
rect 239944 176745 239979 176773
rect 240007 176745 240041 176773
rect 240069 176745 240104 176773
rect 239944 176728 240104 176745
rect 32584 173959 32744 173976
rect 32584 173931 32619 173959
rect 32647 173931 32681 173959
rect 32709 173931 32744 173959
rect 32584 173897 32744 173931
rect 32584 173869 32619 173897
rect 32647 173869 32681 173897
rect 32709 173869 32744 173897
rect 32584 173835 32744 173869
rect 32584 173807 32619 173835
rect 32647 173807 32681 173835
rect 32709 173807 32744 173835
rect 32584 173773 32744 173807
rect 32584 173745 32619 173773
rect 32647 173745 32681 173773
rect 32709 173745 32744 173773
rect 32584 173728 32744 173745
rect 47944 173959 48104 173976
rect 47944 173931 47979 173959
rect 48007 173931 48041 173959
rect 48069 173931 48104 173959
rect 47944 173897 48104 173931
rect 47944 173869 47979 173897
rect 48007 173869 48041 173897
rect 48069 173869 48104 173897
rect 47944 173835 48104 173869
rect 47944 173807 47979 173835
rect 48007 173807 48041 173835
rect 48069 173807 48104 173835
rect 47944 173773 48104 173807
rect 47944 173745 47979 173773
rect 48007 173745 48041 173773
rect 48069 173745 48104 173773
rect 47944 173728 48104 173745
rect 63304 173959 63464 173976
rect 63304 173931 63339 173959
rect 63367 173931 63401 173959
rect 63429 173931 63464 173959
rect 63304 173897 63464 173931
rect 63304 173869 63339 173897
rect 63367 173869 63401 173897
rect 63429 173869 63464 173897
rect 63304 173835 63464 173869
rect 63304 173807 63339 173835
rect 63367 173807 63401 173835
rect 63429 173807 63464 173835
rect 63304 173773 63464 173807
rect 63304 173745 63339 173773
rect 63367 173745 63401 173773
rect 63429 173745 63464 173773
rect 63304 173728 63464 173745
rect 78664 173959 78824 173976
rect 78664 173931 78699 173959
rect 78727 173931 78761 173959
rect 78789 173931 78824 173959
rect 78664 173897 78824 173931
rect 78664 173869 78699 173897
rect 78727 173869 78761 173897
rect 78789 173869 78824 173897
rect 78664 173835 78824 173869
rect 78664 173807 78699 173835
rect 78727 173807 78761 173835
rect 78789 173807 78824 173835
rect 78664 173773 78824 173807
rect 78664 173745 78699 173773
rect 78727 173745 78761 173773
rect 78789 173745 78824 173773
rect 78664 173728 78824 173745
rect 94024 173959 94184 173976
rect 94024 173931 94059 173959
rect 94087 173931 94121 173959
rect 94149 173931 94184 173959
rect 94024 173897 94184 173931
rect 94024 173869 94059 173897
rect 94087 173869 94121 173897
rect 94149 173869 94184 173897
rect 94024 173835 94184 173869
rect 94024 173807 94059 173835
rect 94087 173807 94121 173835
rect 94149 173807 94184 173835
rect 94024 173773 94184 173807
rect 94024 173745 94059 173773
rect 94087 173745 94121 173773
rect 94149 173745 94184 173773
rect 94024 173728 94184 173745
rect 109384 173959 109544 173976
rect 109384 173931 109419 173959
rect 109447 173931 109481 173959
rect 109509 173931 109544 173959
rect 109384 173897 109544 173931
rect 109384 173869 109419 173897
rect 109447 173869 109481 173897
rect 109509 173869 109544 173897
rect 109384 173835 109544 173869
rect 109384 173807 109419 173835
rect 109447 173807 109481 173835
rect 109509 173807 109544 173835
rect 109384 173773 109544 173807
rect 109384 173745 109419 173773
rect 109447 173745 109481 173773
rect 109509 173745 109544 173773
rect 109384 173728 109544 173745
rect 124744 173959 124904 173976
rect 124744 173931 124779 173959
rect 124807 173931 124841 173959
rect 124869 173931 124904 173959
rect 124744 173897 124904 173931
rect 124744 173869 124779 173897
rect 124807 173869 124841 173897
rect 124869 173869 124904 173897
rect 124744 173835 124904 173869
rect 124744 173807 124779 173835
rect 124807 173807 124841 173835
rect 124869 173807 124904 173835
rect 124744 173773 124904 173807
rect 124744 173745 124779 173773
rect 124807 173745 124841 173773
rect 124869 173745 124904 173773
rect 124744 173728 124904 173745
rect 140104 173959 140264 173976
rect 140104 173931 140139 173959
rect 140167 173931 140201 173959
rect 140229 173931 140264 173959
rect 140104 173897 140264 173931
rect 140104 173869 140139 173897
rect 140167 173869 140201 173897
rect 140229 173869 140264 173897
rect 140104 173835 140264 173869
rect 140104 173807 140139 173835
rect 140167 173807 140201 173835
rect 140229 173807 140264 173835
rect 140104 173773 140264 173807
rect 140104 173745 140139 173773
rect 140167 173745 140201 173773
rect 140229 173745 140264 173773
rect 140104 173728 140264 173745
rect 155464 173959 155624 173976
rect 155464 173931 155499 173959
rect 155527 173931 155561 173959
rect 155589 173931 155624 173959
rect 155464 173897 155624 173931
rect 155464 173869 155499 173897
rect 155527 173869 155561 173897
rect 155589 173869 155624 173897
rect 155464 173835 155624 173869
rect 155464 173807 155499 173835
rect 155527 173807 155561 173835
rect 155589 173807 155624 173835
rect 155464 173773 155624 173807
rect 155464 173745 155499 173773
rect 155527 173745 155561 173773
rect 155589 173745 155624 173773
rect 155464 173728 155624 173745
rect 170824 173959 170984 173976
rect 170824 173931 170859 173959
rect 170887 173931 170921 173959
rect 170949 173931 170984 173959
rect 170824 173897 170984 173931
rect 170824 173869 170859 173897
rect 170887 173869 170921 173897
rect 170949 173869 170984 173897
rect 170824 173835 170984 173869
rect 170824 173807 170859 173835
rect 170887 173807 170921 173835
rect 170949 173807 170984 173835
rect 170824 173773 170984 173807
rect 170824 173745 170859 173773
rect 170887 173745 170921 173773
rect 170949 173745 170984 173773
rect 170824 173728 170984 173745
rect 186184 173959 186344 173976
rect 186184 173931 186219 173959
rect 186247 173931 186281 173959
rect 186309 173931 186344 173959
rect 186184 173897 186344 173931
rect 186184 173869 186219 173897
rect 186247 173869 186281 173897
rect 186309 173869 186344 173897
rect 186184 173835 186344 173869
rect 186184 173807 186219 173835
rect 186247 173807 186281 173835
rect 186309 173807 186344 173835
rect 186184 173773 186344 173807
rect 186184 173745 186219 173773
rect 186247 173745 186281 173773
rect 186309 173745 186344 173773
rect 186184 173728 186344 173745
rect 201544 173959 201704 173976
rect 201544 173931 201579 173959
rect 201607 173931 201641 173959
rect 201669 173931 201704 173959
rect 201544 173897 201704 173931
rect 201544 173869 201579 173897
rect 201607 173869 201641 173897
rect 201669 173869 201704 173897
rect 201544 173835 201704 173869
rect 201544 173807 201579 173835
rect 201607 173807 201641 173835
rect 201669 173807 201704 173835
rect 201544 173773 201704 173807
rect 201544 173745 201579 173773
rect 201607 173745 201641 173773
rect 201669 173745 201704 173773
rect 201544 173728 201704 173745
rect 216904 173959 217064 173976
rect 216904 173931 216939 173959
rect 216967 173931 217001 173959
rect 217029 173931 217064 173959
rect 216904 173897 217064 173931
rect 216904 173869 216939 173897
rect 216967 173869 217001 173897
rect 217029 173869 217064 173897
rect 216904 173835 217064 173869
rect 216904 173807 216939 173835
rect 216967 173807 217001 173835
rect 217029 173807 217064 173835
rect 216904 173773 217064 173807
rect 216904 173745 216939 173773
rect 216967 173745 217001 173773
rect 217029 173745 217064 173773
rect 216904 173728 217064 173745
rect 232264 173959 232424 173976
rect 232264 173931 232299 173959
rect 232327 173931 232361 173959
rect 232389 173931 232424 173959
rect 232264 173897 232424 173931
rect 232264 173869 232299 173897
rect 232327 173869 232361 173897
rect 232389 173869 232424 173897
rect 232264 173835 232424 173869
rect 232264 173807 232299 173835
rect 232327 173807 232361 173835
rect 232389 173807 232424 173835
rect 232264 173773 232424 173807
rect 232264 173745 232299 173773
rect 232327 173745 232361 173773
rect 232389 173745 232424 173773
rect 232264 173728 232424 173745
rect 247624 173959 247784 173976
rect 247624 173931 247659 173959
rect 247687 173931 247721 173959
rect 247749 173931 247784 173959
rect 247624 173897 247784 173931
rect 247624 173869 247659 173897
rect 247687 173869 247721 173897
rect 247749 173869 247784 173897
rect 247624 173835 247784 173869
rect 247624 173807 247659 173835
rect 247687 173807 247721 173835
rect 247749 173807 247784 173835
rect 247624 173773 247784 173807
rect 247624 173745 247659 173773
rect 247687 173745 247721 173773
rect 247749 173745 247784 173773
rect 247624 173728 247784 173745
rect 254529 173959 254839 182745
rect 254529 173931 254577 173959
rect 254605 173931 254639 173959
rect 254667 173931 254701 173959
rect 254729 173931 254763 173959
rect 254791 173931 254839 173959
rect 254529 173897 254839 173931
rect 254529 173869 254577 173897
rect 254605 173869 254639 173897
rect 254667 173869 254701 173897
rect 254729 173869 254763 173897
rect 254791 173869 254839 173897
rect 254529 173835 254839 173869
rect 254529 173807 254577 173835
rect 254605 173807 254639 173835
rect 254667 173807 254701 173835
rect 254729 173807 254763 173835
rect 254791 173807 254839 173835
rect 254529 173773 254839 173807
rect 254529 173745 254577 173773
rect 254605 173745 254639 173773
rect 254667 173745 254701 173773
rect 254729 173745 254763 173773
rect 254791 173745 254839 173773
rect 31389 167931 31437 167959
rect 31465 167931 31499 167959
rect 31527 167931 31561 167959
rect 31589 167931 31623 167959
rect 31651 167931 31699 167959
rect 31389 167897 31699 167931
rect 31389 167869 31437 167897
rect 31465 167869 31499 167897
rect 31527 167869 31561 167897
rect 31589 167869 31623 167897
rect 31651 167869 31699 167897
rect 31389 167835 31699 167869
rect 31389 167807 31437 167835
rect 31465 167807 31499 167835
rect 31527 167807 31561 167835
rect 31589 167807 31623 167835
rect 31651 167807 31699 167835
rect 31389 167773 31699 167807
rect 31389 167745 31437 167773
rect 31465 167745 31499 167773
rect 31527 167745 31561 167773
rect 31589 167745 31623 167773
rect 31651 167745 31699 167773
rect 31389 158959 31699 167745
rect 40264 167959 40424 167976
rect 40264 167931 40299 167959
rect 40327 167931 40361 167959
rect 40389 167931 40424 167959
rect 40264 167897 40424 167931
rect 40264 167869 40299 167897
rect 40327 167869 40361 167897
rect 40389 167869 40424 167897
rect 40264 167835 40424 167869
rect 40264 167807 40299 167835
rect 40327 167807 40361 167835
rect 40389 167807 40424 167835
rect 40264 167773 40424 167807
rect 40264 167745 40299 167773
rect 40327 167745 40361 167773
rect 40389 167745 40424 167773
rect 40264 167728 40424 167745
rect 55624 167959 55784 167976
rect 55624 167931 55659 167959
rect 55687 167931 55721 167959
rect 55749 167931 55784 167959
rect 55624 167897 55784 167931
rect 55624 167869 55659 167897
rect 55687 167869 55721 167897
rect 55749 167869 55784 167897
rect 55624 167835 55784 167869
rect 55624 167807 55659 167835
rect 55687 167807 55721 167835
rect 55749 167807 55784 167835
rect 55624 167773 55784 167807
rect 55624 167745 55659 167773
rect 55687 167745 55721 167773
rect 55749 167745 55784 167773
rect 55624 167728 55784 167745
rect 70984 167959 71144 167976
rect 70984 167931 71019 167959
rect 71047 167931 71081 167959
rect 71109 167931 71144 167959
rect 70984 167897 71144 167931
rect 70984 167869 71019 167897
rect 71047 167869 71081 167897
rect 71109 167869 71144 167897
rect 70984 167835 71144 167869
rect 70984 167807 71019 167835
rect 71047 167807 71081 167835
rect 71109 167807 71144 167835
rect 70984 167773 71144 167807
rect 70984 167745 71019 167773
rect 71047 167745 71081 167773
rect 71109 167745 71144 167773
rect 70984 167728 71144 167745
rect 86344 167959 86504 167976
rect 86344 167931 86379 167959
rect 86407 167931 86441 167959
rect 86469 167931 86504 167959
rect 86344 167897 86504 167931
rect 86344 167869 86379 167897
rect 86407 167869 86441 167897
rect 86469 167869 86504 167897
rect 86344 167835 86504 167869
rect 86344 167807 86379 167835
rect 86407 167807 86441 167835
rect 86469 167807 86504 167835
rect 86344 167773 86504 167807
rect 86344 167745 86379 167773
rect 86407 167745 86441 167773
rect 86469 167745 86504 167773
rect 86344 167728 86504 167745
rect 101704 167959 101864 167976
rect 101704 167931 101739 167959
rect 101767 167931 101801 167959
rect 101829 167931 101864 167959
rect 101704 167897 101864 167931
rect 101704 167869 101739 167897
rect 101767 167869 101801 167897
rect 101829 167869 101864 167897
rect 101704 167835 101864 167869
rect 101704 167807 101739 167835
rect 101767 167807 101801 167835
rect 101829 167807 101864 167835
rect 101704 167773 101864 167807
rect 101704 167745 101739 167773
rect 101767 167745 101801 167773
rect 101829 167745 101864 167773
rect 101704 167728 101864 167745
rect 117064 167959 117224 167976
rect 117064 167931 117099 167959
rect 117127 167931 117161 167959
rect 117189 167931 117224 167959
rect 117064 167897 117224 167931
rect 117064 167869 117099 167897
rect 117127 167869 117161 167897
rect 117189 167869 117224 167897
rect 117064 167835 117224 167869
rect 117064 167807 117099 167835
rect 117127 167807 117161 167835
rect 117189 167807 117224 167835
rect 117064 167773 117224 167807
rect 117064 167745 117099 167773
rect 117127 167745 117161 167773
rect 117189 167745 117224 167773
rect 117064 167728 117224 167745
rect 132424 167959 132584 167976
rect 132424 167931 132459 167959
rect 132487 167931 132521 167959
rect 132549 167931 132584 167959
rect 132424 167897 132584 167931
rect 132424 167869 132459 167897
rect 132487 167869 132521 167897
rect 132549 167869 132584 167897
rect 132424 167835 132584 167869
rect 132424 167807 132459 167835
rect 132487 167807 132521 167835
rect 132549 167807 132584 167835
rect 132424 167773 132584 167807
rect 132424 167745 132459 167773
rect 132487 167745 132521 167773
rect 132549 167745 132584 167773
rect 132424 167728 132584 167745
rect 147784 167959 147944 167976
rect 147784 167931 147819 167959
rect 147847 167931 147881 167959
rect 147909 167931 147944 167959
rect 147784 167897 147944 167931
rect 147784 167869 147819 167897
rect 147847 167869 147881 167897
rect 147909 167869 147944 167897
rect 147784 167835 147944 167869
rect 147784 167807 147819 167835
rect 147847 167807 147881 167835
rect 147909 167807 147944 167835
rect 147784 167773 147944 167807
rect 147784 167745 147819 167773
rect 147847 167745 147881 167773
rect 147909 167745 147944 167773
rect 147784 167728 147944 167745
rect 163144 167959 163304 167976
rect 163144 167931 163179 167959
rect 163207 167931 163241 167959
rect 163269 167931 163304 167959
rect 163144 167897 163304 167931
rect 163144 167869 163179 167897
rect 163207 167869 163241 167897
rect 163269 167869 163304 167897
rect 163144 167835 163304 167869
rect 163144 167807 163179 167835
rect 163207 167807 163241 167835
rect 163269 167807 163304 167835
rect 163144 167773 163304 167807
rect 163144 167745 163179 167773
rect 163207 167745 163241 167773
rect 163269 167745 163304 167773
rect 163144 167728 163304 167745
rect 178504 167959 178664 167976
rect 178504 167931 178539 167959
rect 178567 167931 178601 167959
rect 178629 167931 178664 167959
rect 178504 167897 178664 167931
rect 178504 167869 178539 167897
rect 178567 167869 178601 167897
rect 178629 167869 178664 167897
rect 178504 167835 178664 167869
rect 178504 167807 178539 167835
rect 178567 167807 178601 167835
rect 178629 167807 178664 167835
rect 178504 167773 178664 167807
rect 178504 167745 178539 167773
rect 178567 167745 178601 167773
rect 178629 167745 178664 167773
rect 178504 167728 178664 167745
rect 193864 167959 194024 167976
rect 193864 167931 193899 167959
rect 193927 167931 193961 167959
rect 193989 167931 194024 167959
rect 193864 167897 194024 167931
rect 193864 167869 193899 167897
rect 193927 167869 193961 167897
rect 193989 167869 194024 167897
rect 193864 167835 194024 167869
rect 193864 167807 193899 167835
rect 193927 167807 193961 167835
rect 193989 167807 194024 167835
rect 193864 167773 194024 167807
rect 193864 167745 193899 167773
rect 193927 167745 193961 167773
rect 193989 167745 194024 167773
rect 193864 167728 194024 167745
rect 209224 167959 209384 167976
rect 209224 167931 209259 167959
rect 209287 167931 209321 167959
rect 209349 167931 209384 167959
rect 209224 167897 209384 167931
rect 209224 167869 209259 167897
rect 209287 167869 209321 167897
rect 209349 167869 209384 167897
rect 209224 167835 209384 167869
rect 209224 167807 209259 167835
rect 209287 167807 209321 167835
rect 209349 167807 209384 167835
rect 209224 167773 209384 167807
rect 209224 167745 209259 167773
rect 209287 167745 209321 167773
rect 209349 167745 209384 167773
rect 209224 167728 209384 167745
rect 224584 167959 224744 167976
rect 224584 167931 224619 167959
rect 224647 167931 224681 167959
rect 224709 167931 224744 167959
rect 224584 167897 224744 167931
rect 224584 167869 224619 167897
rect 224647 167869 224681 167897
rect 224709 167869 224744 167897
rect 224584 167835 224744 167869
rect 224584 167807 224619 167835
rect 224647 167807 224681 167835
rect 224709 167807 224744 167835
rect 224584 167773 224744 167807
rect 224584 167745 224619 167773
rect 224647 167745 224681 167773
rect 224709 167745 224744 167773
rect 224584 167728 224744 167745
rect 239944 167959 240104 167976
rect 239944 167931 239979 167959
rect 240007 167931 240041 167959
rect 240069 167931 240104 167959
rect 239944 167897 240104 167931
rect 239944 167869 239979 167897
rect 240007 167869 240041 167897
rect 240069 167869 240104 167897
rect 239944 167835 240104 167869
rect 239944 167807 239979 167835
rect 240007 167807 240041 167835
rect 240069 167807 240104 167835
rect 239944 167773 240104 167807
rect 239944 167745 239979 167773
rect 240007 167745 240041 167773
rect 240069 167745 240104 167773
rect 239944 167728 240104 167745
rect 32584 164959 32744 164976
rect 32584 164931 32619 164959
rect 32647 164931 32681 164959
rect 32709 164931 32744 164959
rect 32584 164897 32744 164931
rect 32584 164869 32619 164897
rect 32647 164869 32681 164897
rect 32709 164869 32744 164897
rect 32584 164835 32744 164869
rect 32584 164807 32619 164835
rect 32647 164807 32681 164835
rect 32709 164807 32744 164835
rect 32584 164773 32744 164807
rect 32584 164745 32619 164773
rect 32647 164745 32681 164773
rect 32709 164745 32744 164773
rect 32584 164728 32744 164745
rect 47944 164959 48104 164976
rect 47944 164931 47979 164959
rect 48007 164931 48041 164959
rect 48069 164931 48104 164959
rect 47944 164897 48104 164931
rect 47944 164869 47979 164897
rect 48007 164869 48041 164897
rect 48069 164869 48104 164897
rect 47944 164835 48104 164869
rect 47944 164807 47979 164835
rect 48007 164807 48041 164835
rect 48069 164807 48104 164835
rect 47944 164773 48104 164807
rect 47944 164745 47979 164773
rect 48007 164745 48041 164773
rect 48069 164745 48104 164773
rect 47944 164728 48104 164745
rect 63304 164959 63464 164976
rect 63304 164931 63339 164959
rect 63367 164931 63401 164959
rect 63429 164931 63464 164959
rect 63304 164897 63464 164931
rect 63304 164869 63339 164897
rect 63367 164869 63401 164897
rect 63429 164869 63464 164897
rect 63304 164835 63464 164869
rect 63304 164807 63339 164835
rect 63367 164807 63401 164835
rect 63429 164807 63464 164835
rect 63304 164773 63464 164807
rect 63304 164745 63339 164773
rect 63367 164745 63401 164773
rect 63429 164745 63464 164773
rect 63304 164728 63464 164745
rect 78664 164959 78824 164976
rect 78664 164931 78699 164959
rect 78727 164931 78761 164959
rect 78789 164931 78824 164959
rect 78664 164897 78824 164931
rect 78664 164869 78699 164897
rect 78727 164869 78761 164897
rect 78789 164869 78824 164897
rect 78664 164835 78824 164869
rect 78664 164807 78699 164835
rect 78727 164807 78761 164835
rect 78789 164807 78824 164835
rect 78664 164773 78824 164807
rect 78664 164745 78699 164773
rect 78727 164745 78761 164773
rect 78789 164745 78824 164773
rect 78664 164728 78824 164745
rect 94024 164959 94184 164976
rect 94024 164931 94059 164959
rect 94087 164931 94121 164959
rect 94149 164931 94184 164959
rect 94024 164897 94184 164931
rect 94024 164869 94059 164897
rect 94087 164869 94121 164897
rect 94149 164869 94184 164897
rect 94024 164835 94184 164869
rect 94024 164807 94059 164835
rect 94087 164807 94121 164835
rect 94149 164807 94184 164835
rect 94024 164773 94184 164807
rect 94024 164745 94059 164773
rect 94087 164745 94121 164773
rect 94149 164745 94184 164773
rect 94024 164728 94184 164745
rect 109384 164959 109544 164976
rect 109384 164931 109419 164959
rect 109447 164931 109481 164959
rect 109509 164931 109544 164959
rect 109384 164897 109544 164931
rect 109384 164869 109419 164897
rect 109447 164869 109481 164897
rect 109509 164869 109544 164897
rect 109384 164835 109544 164869
rect 109384 164807 109419 164835
rect 109447 164807 109481 164835
rect 109509 164807 109544 164835
rect 109384 164773 109544 164807
rect 109384 164745 109419 164773
rect 109447 164745 109481 164773
rect 109509 164745 109544 164773
rect 109384 164728 109544 164745
rect 124744 164959 124904 164976
rect 124744 164931 124779 164959
rect 124807 164931 124841 164959
rect 124869 164931 124904 164959
rect 124744 164897 124904 164931
rect 124744 164869 124779 164897
rect 124807 164869 124841 164897
rect 124869 164869 124904 164897
rect 124744 164835 124904 164869
rect 124744 164807 124779 164835
rect 124807 164807 124841 164835
rect 124869 164807 124904 164835
rect 124744 164773 124904 164807
rect 124744 164745 124779 164773
rect 124807 164745 124841 164773
rect 124869 164745 124904 164773
rect 124744 164728 124904 164745
rect 140104 164959 140264 164976
rect 140104 164931 140139 164959
rect 140167 164931 140201 164959
rect 140229 164931 140264 164959
rect 140104 164897 140264 164931
rect 140104 164869 140139 164897
rect 140167 164869 140201 164897
rect 140229 164869 140264 164897
rect 140104 164835 140264 164869
rect 140104 164807 140139 164835
rect 140167 164807 140201 164835
rect 140229 164807 140264 164835
rect 140104 164773 140264 164807
rect 140104 164745 140139 164773
rect 140167 164745 140201 164773
rect 140229 164745 140264 164773
rect 140104 164728 140264 164745
rect 155464 164959 155624 164976
rect 155464 164931 155499 164959
rect 155527 164931 155561 164959
rect 155589 164931 155624 164959
rect 155464 164897 155624 164931
rect 155464 164869 155499 164897
rect 155527 164869 155561 164897
rect 155589 164869 155624 164897
rect 155464 164835 155624 164869
rect 155464 164807 155499 164835
rect 155527 164807 155561 164835
rect 155589 164807 155624 164835
rect 155464 164773 155624 164807
rect 155464 164745 155499 164773
rect 155527 164745 155561 164773
rect 155589 164745 155624 164773
rect 155464 164728 155624 164745
rect 170824 164959 170984 164976
rect 170824 164931 170859 164959
rect 170887 164931 170921 164959
rect 170949 164931 170984 164959
rect 170824 164897 170984 164931
rect 170824 164869 170859 164897
rect 170887 164869 170921 164897
rect 170949 164869 170984 164897
rect 170824 164835 170984 164869
rect 170824 164807 170859 164835
rect 170887 164807 170921 164835
rect 170949 164807 170984 164835
rect 170824 164773 170984 164807
rect 170824 164745 170859 164773
rect 170887 164745 170921 164773
rect 170949 164745 170984 164773
rect 170824 164728 170984 164745
rect 186184 164959 186344 164976
rect 186184 164931 186219 164959
rect 186247 164931 186281 164959
rect 186309 164931 186344 164959
rect 186184 164897 186344 164931
rect 186184 164869 186219 164897
rect 186247 164869 186281 164897
rect 186309 164869 186344 164897
rect 186184 164835 186344 164869
rect 186184 164807 186219 164835
rect 186247 164807 186281 164835
rect 186309 164807 186344 164835
rect 186184 164773 186344 164807
rect 186184 164745 186219 164773
rect 186247 164745 186281 164773
rect 186309 164745 186344 164773
rect 186184 164728 186344 164745
rect 201544 164959 201704 164976
rect 201544 164931 201579 164959
rect 201607 164931 201641 164959
rect 201669 164931 201704 164959
rect 201544 164897 201704 164931
rect 201544 164869 201579 164897
rect 201607 164869 201641 164897
rect 201669 164869 201704 164897
rect 201544 164835 201704 164869
rect 201544 164807 201579 164835
rect 201607 164807 201641 164835
rect 201669 164807 201704 164835
rect 201544 164773 201704 164807
rect 201544 164745 201579 164773
rect 201607 164745 201641 164773
rect 201669 164745 201704 164773
rect 201544 164728 201704 164745
rect 216904 164959 217064 164976
rect 216904 164931 216939 164959
rect 216967 164931 217001 164959
rect 217029 164931 217064 164959
rect 216904 164897 217064 164931
rect 216904 164869 216939 164897
rect 216967 164869 217001 164897
rect 217029 164869 217064 164897
rect 216904 164835 217064 164869
rect 216904 164807 216939 164835
rect 216967 164807 217001 164835
rect 217029 164807 217064 164835
rect 216904 164773 217064 164807
rect 216904 164745 216939 164773
rect 216967 164745 217001 164773
rect 217029 164745 217064 164773
rect 216904 164728 217064 164745
rect 232264 164959 232424 164976
rect 232264 164931 232299 164959
rect 232327 164931 232361 164959
rect 232389 164931 232424 164959
rect 232264 164897 232424 164931
rect 232264 164869 232299 164897
rect 232327 164869 232361 164897
rect 232389 164869 232424 164897
rect 232264 164835 232424 164869
rect 232264 164807 232299 164835
rect 232327 164807 232361 164835
rect 232389 164807 232424 164835
rect 232264 164773 232424 164807
rect 232264 164745 232299 164773
rect 232327 164745 232361 164773
rect 232389 164745 232424 164773
rect 232264 164728 232424 164745
rect 247624 164959 247784 164976
rect 247624 164931 247659 164959
rect 247687 164931 247721 164959
rect 247749 164931 247784 164959
rect 247624 164897 247784 164931
rect 247624 164869 247659 164897
rect 247687 164869 247721 164897
rect 247749 164869 247784 164897
rect 247624 164835 247784 164869
rect 247624 164807 247659 164835
rect 247687 164807 247721 164835
rect 247749 164807 247784 164835
rect 247624 164773 247784 164807
rect 247624 164745 247659 164773
rect 247687 164745 247721 164773
rect 247749 164745 247784 164773
rect 247624 164728 247784 164745
rect 254529 164959 254839 173745
rect 254529 164931 254577 164959
rect 254605 164931 254639 164959
rect 254667 164931 254701 164959
rect 254729 164931 254763 164959
rect 254791 164931 254839 164959
rect 254529 164897 254839 164931
rect 254529 164869 254577 164897
rect 254605 164869 254639 164897
rect 254667 164869 254701 164897
rect 254729 164869 254763 164897
rect 254791 164869 254839 164897
rect 254529 164835 254839 164869
rect 254529 164807 254577 164835
rect 254605 164807 254639 164835
rect 254667 164807 254701 164835
rect 254729 164807 254763 164835
rect 254791 164807 254839 164835
rect 254529 164773 254839 164807
rect 254529 164745 254577 164773
rect 254605 164745 254639 164773
rect 254667 164745 254701 164773
rect 254729 164745 254763 164773
rect 254791 164745 254839 164773
rect 31389 158931 31437 158959
rect 31465 158931 31499 158959
rect 31527 158931 31561 158959
rect 31589 158931 31623 158959
rect 31651 158931 31699 158959
rect 31389 158897 31699 158931
rect 31389 158869 31437 158897
rect 31465 158869 31499 158897
rect 31527 158869 31561 158897
rect 31589 158869 31623 158897
rect 31651 158869 31699 158897
rect 31389 158835 31699 158869
rect 31389 158807 31437 158835
rect 31465 158807 31499 158835
rect 31527 158807 31561 158835
rect 31589 158807 31623 158835
rect 31651 158807 31699 158835
rect 31389 158773 31699 158807
rect 31389 158745 31437 158773
rect 31465 158745 31499 158773
rect 31527 158745 31561 158773
rect 31589 158745 31623 158773
rect 31651 158745 31699 158773
rect 31389 149959 31699 158745
rect 40264 158959 40424 158976
rect 40264 158931 40299 158959
rect 40327 158931 40361 158959
rect 40389 158931 40424 158959
rect 40264 158897 40424 158931
rect 40264 158869 40299 158897
rect 40327 158869 40361 158897
rect 40389 158869 40424 158897
rect 40264 158835 40424 158869
rect 40264 158807 40299 158835
rect 40327 158807 40361 158835
rect 40389 158807 40424 158835
rect 40264 158773 40424 158807
rect 40264 158745 40299 158773
rect 40327 158745 40361 158773
rect 40389 158745 40424 158773
rect 40264 158728 40424 158745
rect 55624 158959 55784 158976
rect 55624 158931 55659 158959
rect 55687 158931 55721 158959
rect 55749 158931 55784 158959
rect 55624 158897 55784 158931
rect 55624 158869 55659 158897
rect 55687 158869 55721 158897
rect 55749 158869 55784 158897
rect 55624 158835 55784 158869
rect 55624 158807 55659 158835
rect 55687 158807 55721 158835
rect 55749 158807 55784 158835
rect 55624 158773 55784 158807
rect 55624 158745 55659 158773
rect 55687 158745 55721 158773
rect 55749 158745 55784 158773
rect 55624 158728 55784 158745
rect 70984 158959 71144 158976
rect 70984 158931 71019 158959
rect 71047 158931 71081 158959
rect 71109 158931 71144 158959
rect 70984 158897 71144 158931
rect 70984 158869 71019 158897
rect 71047 158869 71081 158897
rect 71109 158869 71144 158897
rect 70984 158835 71144 158869
rect 70984 158807 71019 158835
rect 71047 158807 71081 158835
rect 71109 158807 71144 158835
rect 70984 158773 71144 158807
rect 70984 158745 71019 158773
rect 71047 158745 71081 158773
rect 71109 158745 71144 158773
rect 70984 158728 71144 158745
rect 86344 158959 86504 158976
rect 86344 158931 86379 158959
rect 86407 158931 86441 158959
rect 86469 158931 86504 158959
rect 86344 158897 86504 158931
rect 86344 158869 86379 158897
rect 86407 158869 86441 158897
rect 86469 158869 86504 158897
rect 86344 158835 86504 158869
rect 86344 158807 86379 158835
rect 86407 158807 86441 158835
rect 86469 158807 86504 158835
rect 86344 158773 86504 158807
rect 86344 158745 86379 158773
rect 86407 158745 86441 158773
rect 86469 158745 86504 158773
rect 86344 158728 86504 158745
rect 101704 158959 101864 158976
rect 101704 158931 101739 158959
rect 101767 158931 101801 158959
rect 101829 158931 101864 158959
rect 101704 158897 101864 158931
rect 101704 158869 101739 158897
rect 101767 158869 101801 158897
rect 101829 158869 101864 158897
rect 101704 158835 101864 158869
rect 101704 158807 101739 158835
rect 101767 158807 101801 158835
rect 101829 158807 101864 158835
rect 101704 158773 101864 158807
rect 101704 158745 101739 158773
rect 101767 158745 101801 158773
rect 101829 158745 101864 158773
rect 101704 158728 101864 158745
rect 117064 158959 117224 158976
rect 117064 158931 117099 158959
rect 117127 158931 117161 158959
rect 117189 158931 117224 158959
rect 117064 158897 117224 158931
rect 117064 158869 117099 158897
rect 117127 158869 117161 158897
rect 117189 158869 117224 158897
rect 117064 158835 117224 158869
rect 117064 158807 117099 158835
rect 117127 158807 117161 158835
rect 117189 158807 117224 158835
rect 117064 158773 117224 158807
rect 117064 158745 117099 158773
rect 117127 158745 117161 158773
rect 117189 158745 117224 158773
rect 117064 158728 117224 158745
rect 132424 158959 132584 158976
rect 132424 158931 132459 158959
rect 132487 158931 132521 158959
rect 132549 158931 132584 158959
rect 132424 158897 132584 158931
rect 132424 158869 132459 158897
rect 132487 158869 132521 158897
rect 132549 158869 132584 158897
rect 132424 158835 132584 158869
rect 132424 158807 132459 158835
rect 132487 158807 132521 158835
rect 132549 158807 132584 158835
rect 132424 158773 132584 158807
rect 132424 158745 132459 158773
rect 132487 158745 132521 158773
rect 132549 158745 132584 158773
rect 132424 158728 132584 158745
rect 147784 158959 147944 158976
rect 147784 158931 147819 158959
rect 147847 158931 147881 158959
rect 147909 158931 147944 158959
rect 147784 158897 147944 158931
rect 147784 158869 147819 158897
rect 147847 158869 147881 158897
rect 147909 158869 147944 158897
rect 147784 158835 147944 158869
rect 147784 158807 147819 158835
rect 147847 158807 147881 158835
rect 147909 158807 147944 158835
rect 147784 158773 147944 158807
rect 147784 158745 147819 158773
rect 147847 158745 147881 158773
rect 147909 158745 147944 158773
rect 147784 158728 147944 158745
rect 163144 158959 163304 158976
rect 163144 158931 163179 158959
rect 163207 158931 163241 158959
rect 163269 158931 163304 158959
rect 163144 158897 163304 158931
rect 163144 158869 163179 158897
rect 163207 158869 163241 158897
rect 163269 158869 163304 158897
rect 163144 158835 163304 158869
rect 163144 158807 163179 158835
rect 163207 158807 163241 158835
rect 163269 158807 163304 158835
rect 163144 158773 163304 158807
rect 163144 158745 163179 158773
rect 163207 158745 163241 158773
rect 163269 158745 163304 158773
rect 163144 158728 163304 158745
rect 178504 158959 178664 158976
rect 178504 158931 178539 158959
rect 178567 158931 178601 158959
rect 178629 158931 178664 158959
rect 178504 158897 178664 158931
rect 178504 158869 178539 158897
rect 178567 158869 178601 158897
rect 178629 158869 178664 158897
rect 178504 158835 178664 158869
rect 178504 158807 178539 158835
rect 178567 158807 178601 158835
rect 178629 158807 178664 158835
rect 178504 158773 178664 158807
rect 178504 158745 178539 158773
rect 178567 158745 178601 158773
rect 178629 158745 178664 158773
rect 178504 158728 178664 158745
rect 193864 158959 194024 158976
rect 193864 158931 193899 158959
rect 193927 158931 193961 158959
rect 193989 158931 194024 158959
rect 193864 158897 194024 158931
rect 193864 158869 193899 158897
rect 193927 158869 193961 158897
rect 193989 158869 194024 158897
rect 193864 158835 194024 158869
rect 193864 158807 193899 158835
rect 193927 158807 193961 158835
rect 193989 158807 194024 158835
rect 193864 158773 194024 158807
rect 193864 158745 193899 158773
rect 193927 158745 193961 158773
rect 193989 158745 194024 158773
rect 193864 158728 194024 158745
rect 209224 158959 209384 158976
rect 209224 158931 209259 158959
rect 209287 158931 209321 158959
rect 209349 158931 209384 158959
rect 209224 158897 209384 158931
rect 209224 158869 209259 158897
rect 209287 158869 209321 158897
rect 209349 158869 209384 158897
rect 209224 158835 209384 158869
rect 209224 158807 209259 158835
rect 209287 158807 209321 158835
rect 209349 158807 209384 158835
rect 209224 158773 209384 158807
rect 209224 158745 209259 158773
rect 209287 158745 209321 158773
rect 209349 158745 209384 158773
rect 209224 158728 209384 158745
rect 224584 158959 224744 158976
rect 224584 158931 224619 158959
rect 224647 158931 224681 158959
rect 224709 158931 224744 158959
rect 224584 158897 224744 158931
rect 224584 158869 224619 158897
rect 224647 158869 224681 158897
rect 224709 158869 224744 158897
rect 224584 158835 224744 158869
rect 224584 158807 224619 158835
rect 224647 158807 224681 158835
rect 224709 158807 224744 158835
rect 224584 158773 224744 158807
rect 224584 158745 224619 158773
rect 224647 158745 224681 158773
rect 224709 158745 224744 158773
rect 224584 158728 224744 158745
rect 239944 158959 240104 158976
rect 239944 158931 239979 158959
rect 240007 158931 240041 158959
rect 240069 158931 240104 158959
rect 239944 158897 240104 158931
rect 239944 158869 239979 158897
rect 240007 158869 240041 158897
rect 240069 158869 240104 158897
rect 239944 158835 240104 158869
rect 239944 158807 239979 158835
rect 240007 158807 240041 158835
rect 240069 158807 240104 158835
rect 239944 158773 240104 158807
rect 239944 158745 239979 158773
rect 240007 158745 240041 158773
rect 240069 158745 240104 158773
rect 239944 158728 240104 158745
rect 32584 155959 32744 155976
rect 32584 155931 32619 155959
rect 32647 155931 32681 155959
rect 32709 155931 32744 155959
rect 32584 155897 32744 155931
rect 32584 155869 32619 155897
rect 32647 155869 32681 155897
rect 32709 155869 32744 155897
rect 32584 155835 32744 155869
rect 32584 155807 32619 155835
rect 32647 155807 32681 155835
rect 32709 155807 32744 155835
rect 32584 155773 32744 155807
rect 32584 155745 32619 155773
rect 32647 155745 32681 155773
rect 32709 155745 32744 155773
rect 32584 155728 32744 155745
rect 47944 155959 48104 155976
rect 47944 155931 47979 155959
rect 48007 155931 48041 155959
rect 48069 155931 48104 155959
rect 47944 155897 48104 155931
rect 47944 155869 47979 155897
rect 48007 155869 48041 155897
rect 48069 155869 48104 155897
rect 47944 155835 48104 155869
rect 47944 155807 47979 155835
rect 48007 155807 48041 155835
rect 48069 155807 48104 155835
rect 47944 155773 48104 155807
rect 47944 155745 47979 155773
rect 48007 155745 48041 155773
rect 48069 155745 48104 155773
rect 47944 155728 48104 155745
rect 63304 155959 63464 155976
rect 63304 155931 63339 155959
rect 63367 155931 63401 155959
rect 63429 155931 63464 155959
rect 63304 155897 63464 155931
rect 63304 155869 63339 155897
rect 63367 155869 63401 155897
rect 63429 155869 63464 155897
rect 63304 155835 63464 155869
rect 63304 155807 63339 155835
rect 63367 155807 63401 155835
rect 63429 155807 63464 155835
rect 63304 155773 63464 155807
rect 63304 155745 63339 155773
rect 63367 155745 63401 155773
rect 63429 155745 63464 155773
rect 63304 155728 63464 155745
rect 78664 155959 78824 155976
rect 78664 155931 78699 155959
rect 78727 155931 78761 155959
rect 78789 155931 78824 155959
rect 78664 155897 78824 155931
rect 78664 155869 78699 155897
rect 78727 155869 78761 155897
rect 78789 155869 78824 155897
rect 78664 155835 78824 155869
rect 78664 155807 78699 155835
rect 78727 155807 78761 155835
rect 78789 155807 78824 155835
rect 78664 155773 78824 155807
rect 78664 155745 78699 155773
rect 78727 155745 78761 155773
rect 78789 155745 78824 155773
rect 78664 155728 78824 155745
rect 94024 155959 94184 155976
rect 94024 155931 94059 155959
rect 94087 155931 94121 155959
rect 94149 155931 94184 155959
rect 94024 155897 94184 155931
rect 94024 155869 94059 155897
rect 94087 155869 94121 155897
rect 94149 155869 94184 155897
rect 94024 155835 94184 155869
rect 94024 155807 94059 155835
rect 94087 155807 94121 155835
rect 94149 155807 94184 155835
rect 94024 155773 94184 155807
rect 94024 155745 94059 155773
rect 94087 155745 94121 155773
rect 94149 155745 94184 155773
rect 94024 155728 94184 155745
rect 109384 155959 109544 155976
rect 109384 155931 109419 155959
rect 109447 155931 109481 155959
rect 109509 155931 109544 155959
rect 109384 155897 109544 155931
rect 109384 155869 109419 155897
rect 109447 155869 109481 155897
rect 109509 155869 109544 155897
rect 109384 155835 109544 155869
rect 109384 155807 109419 155835
rect 109447 155807 109481 155835
rect 109509 155807 109544 155835
rect 109384 155773 109544 155807
rect 109384 155745 109419 155773
rect 109447 155745 109481 155773
rect 109509 155745 109544 155773
rect 109384 155728 109544 155745
rect 124744 155959 124904 155976
rect 124744 155931 124779 155959
rect 124807 155931 124841 155959
rect 124869 155931 124904 155959
rect 124744 155897 124904 155931
rect 124744 155869 124779 155897
rect 124807 155869 124841 155897
rect 124869 155869 124904 155897
rect 124744 155835 124904 155869
rect 124744 155807 124779 155835
rect 124807 155807 124841 155835
rect 124869 155807 124904 155835
rect 124744 155773 124904 155807
rect 124744 155745 124779 155773
rect 124807 155745 124841 155773
rect 124869 155745 124904 155773
rect 124744 155728 124904 155745
rect 140104 155959 140264 155976
rect 140104 155931 140139 155959
rect 140167 155931 140201 155959
rect 140229 155931 140264 155959
rect 140104 155897 140264 155931
rect 140104 155869 140139 155897
rect 140167 155869 140201 155897
rect 140229 155869 140264 155897
rect 140104 155835 140264 155869
rect 140104 155807 140139 155835
rect 140167 155807 140201 155835
rect 140229 155807 140264 155835
rect 140104 155773 140264 155807
rect 140104 155745 140139 155773
rect 140167 155745 140201 155773
rect 140229 155745 140264 155773
rect 140104 155728 140264 155745
rect 155464 155959 155624 155976
rect 155464 155931 155499 155959
rect 155527 155931 155561 155959
rect 155589 155931 155624 155959
rect 155464 155897 155624 155931
rect 155464 155869 155499 155897
rect 155527 155869 155561 155897
rect 155589 155869 155624 155897
rect 155464 155835 155624 155869
rect 155464 155807 155499 155835
rect 155527 155807 155561 155835
rect 155589 155807 155624 155835
rect 155464 155773 155624 155807
rect 155464 155745 155499 155773
rect 155527 155745 155561 155773
rect 155589 155745 155624 155773
rect 155464 155728 155624 155745
rect 170824 155959 170984 155976
rect 170824 155931 170859 155959
rect 170887 155931 170921 155959
rect 170949 155931 170984 155959
rect 170824 155897 170984 155931
rect 170824 155869 170859 155897
rect 170887 155869 170921 155897
rect 170949 155869 170984 155897
rect 170824 155835 170984 155869
rect 170824 155807 170859 155835
rect 170887 155807 170921 155835
rect 170949 155807 170984 155835
rect 170824 155773 170984 155807
rect 170824 155745 170859 155773
rect 170887 155745 170921 155773
rect 170949 155745 170984 155773
rect 170824 155728 170984 155745
rect 186184 155959 186344 155976
rect 186184 155931 186219 155959
rect 186247 155931 186281 155959
rect 186309 155931 186344 155959
rect 186184 155897 186344 155931
rect 186184 155869 186219 155897
rect 186247 155869 186281 155897
rect 186309 155869 186344 155897
rect 186184 155835 186344 155869
rect 186184 155807 186219 155835
rect 186247 155807 186281 155835
rect 186309 155807 186344 155835
rect 186184 155773 186344 155807
rect 186184 155745 186219 155773
rect 186247 155745 186281 155773
rect 186309 155745 186344 155773
rect 186184 155728 186344 155745
rect 201544 155959 201704 155976
rect 201544 155931 201579 155959
rect 201607 155931 201641 155959
rect 201669 155931 201704 155959
rect 201544 155897 201704 155931
rect 201544 155869 201579 155897
rect 201607 155869 201641 155897
rect 201669 155869 201704 155897
rect 201544 155835 201704 155869
rect 201544 155807 201579 155835
rect 201607 155807 201641 155835
rect 201669 155807 201704 155835
rect 201544 155773 201704 155807
rect 201544 155745 201579 155773
rect 201607 155745 201641 155773
rect 201669 155745 201704 155773
rect 201544 155728 201704 155745
rect 216904 155959 217064 155976
rect 216904 155931 216939 155959
rect 216967 155931 217001 155959
rect 217029 155931 217064 155959
rect 216904 155897 217064 155931
rect 216904 155869 216939 155897
rect 216967 155869 217001 155897
rect 217029 155869 217064 155897
rect 216904 155835 217064 155869
rect 216904 155807 216939 155835
rect 216967 155807 217001 155835
rect 217029 155807 217064 155835
rect 216904 155773 217064 155807
rect 216904 155745 216939 155773
rect 216967 155745 217001 155773
rect 217029 155745 217064 155773
rect 216904 155728 217064 155745
rect 232264 155959 232424 155976
rect 232264 155931 232299 155959
rect 232327 155931 232361 155959
rect 232389 155931 232424 155959
rect 232264 155897 232424 155931
rect 232264 155869 232299 155897
rect 232327 155869 232361 155897
rect 232389 155869 232424 155897
rect 232264 155835 232424 155869
rect 232264 155807 232299 155835
rect 232327 155807 232361 155835
rect 232389 155807 232424 155835
rect 232264 155773 232424 155807
rect 232264 155745 232299 155773
rect 232327 155745 232361 155773
rect 232389 155745 232424 155773
rect 232264 155728 232424 155745
rect 247624 155959 247784 155976
rect 247624 155931 247659 155959
rect 247687 155931 247721 155959
rect 247749 155931 247784 155959
rect 247624 155897 247784 155931
rect 247624 155869 247659 155897
rect 247687 155869 247721 155897
rect 247749 155869 247784 155897
rect 247624 155835 247784 155869
rect 247624 155807 247659 155835
rect 247687 155807 247721 155835
rect 247749 155807 247784 155835
rect 247624 155773 247784 155807
rect 247624 155745 247659 155773
rect 247687 155745 247721 155773
rect 247749 155745 247784 155773
rect 247624 155728 247784 155745
rect 254529 155959 254839 164745
rect 254529 155931 254577 155959
rect 254605 155931 254639 155959
rect 254667 155931 254701 155959
rect 254729 155931 254763 155959
rect 254791 155931 254839 155959
rect 254529 155897 254839 155931
rect 254529 155869 254577 155897
rect 254605 155869 254639 155897
rect 254667 155869 254701 155897
rect 254729 155869 254763 155897
rect 254791 155869 254839 155897
rect 254529 155835 254839 155869
rect 254529 155807 254577 155835
rect 254605 155807 254639 155835
rect 254667 155807 254701 155835
rect 254729 155807 254763 155835
rect 254791 155807 254839 155835
rect 254529 155773 254839 155807
rect 254529 155745 254577 155773
rect 254605 155745 254639 155773
rect 254667 155745 254701 155773
rect 254729 155745 254763 155773
rect 254791 155745 254839 155773
rect 31389 149931 31437 149959
rect 31465 149931 31499 149959
rect 31527 149931 31561 149959
rect 31589 149931 31623 149959
rect 31651 149931 31699 149959
rect 31389 149897 31699 149931
rect 31389 149869 31437 149897
rect 31465 149869 31499 149897
rect 31527 149869 31561 149897
rect 31589 149869 31623 149897
rect 31651 149869 31699 149897
rect 31389 149835 31699 149869
rect 31389 149807 31437 149835
rect 31465 149807 31499 149835
rect 31527 149807 31561 149835
rect 31589 149807 31623 149835
rect 31651 149807 31699 149835
rect 31389 149773 31699 149807
rect 31389 149745 31437 149773
rect 31465 149745 31499 149773
rect 31527 149745 31561 149773
rect 31589 149745 31623 149773
rect 31651 149745 31699 149773
rect 31389 140959 31699 149745
rect 40264 149959 40424 149976
rect 40264 149931 40299 149959
rect 40327 149931 40361 149959
rect 40389 149931 40424 149959
rect 40264 149897 40424 149931
rect 40264 149869 40299 149897
rect 40327 149869 40361 149897
rect 40389 149869 40424 149897
rect 40264 149835 40424 149869
rect 40264 149807 40299 149835
rect 40327 149807 40361 149835
rect 40389 149807 40424 149835
rect 40264 149773 40424 149807
rect 40264 149745 40299 149773
rect 40327 149745 40361 149773
rect 40389 149745 40424 149773
rect 40264 149728 40424 149745
rect 55624 149959 55784 149976
rect 55624 149931 55659 149959
rect 55687 149931 55721 149959
rect 55749 149931 55784 149959
rect 55624 149897 55784 149931
rect 55624 149869 55659 149897
rect 55687 149869 55721 149897
rect 55749 149869 55784 149897
rect 55624 149835 55784 149869
rect 55624 149807 55659 149835
rect 55687 149807 55721 149835
rect 55749 149807 55784 149835
rect 55624 149773 55784 149807
rect 55624 149745 55659 149773
rect 55687 149745 55721 149773
rect 55749 149745 55784 149773
rect 55624 149728 55784 149745
rect 70984 149959 71144 149976
rect 70984 149931 71019 149959
rect 71047 149931 71081 149959
rect 71109 149931 71144 149959
rect 70984 149897 71144 149931
rect 70984 149869 71019 149897
rect 71047 149869 71081 149897
rect 71109 149869 71144 149897
rect 70984 149835 71144 149869
rect 70984 149807 71019 149835
rect 71047 149807 71081 149835
rect 71109 149807 71144 149835
rect 70984 149773 71144 149807
rect 70984 149745 71019 149773
rect 71047 149745 71081 149773
rect 71109 149745 71144 149773
rect 70984 149728 71144 149745
rect 86344 149959 86504 149976
rect 86344 149931 86379 149959
rect 86407 149931 86441 149959
rect 86469 149931 86504 149959
rect 86344 149897 86504 149931
rect 86344 149869 86379 149897
rect 86407 149869 86441 149897
rect 86469 149869 86504 149897
rect 86344 149835 86504 149869
rect 86344 149807 86379 149835
rect 86407 149807 86441 149835
rect 86469 149807 86504 149835
rect 86344 149773 86504 149807
rect 86344 149745 86379 149773
rect 86407 149745 86441 149773
rect 86469 149745 86504 149773
rect 86344 149728 86504 149745
rect 101704 149959 101864 149976
rect 101704 149931 101739 149959
rect 101767 149931 101801 149959
rect 101829 149931 101864 149959
rect 101704 149897 101864 149931
rect 101704 149869 101739 149897
rect 101767 149869 101801 149897
rect 101829 149869 101864 149897
rect 101704 149835 101864 149869
rect 101704 149807 101739 149835
rect 101767 149807 101801 149835
rect 101829 149807 101864 149835
rect 101704 149773 101864 149807
rect 101704 149745 101739 149773
rect 101767 149745 101801 149773
rect 101829 149745 101864 149773
rect 101704 149728 101864 149745
rect 117064 149959 117224 149976
rect 117064 149931 117099 149959
rect 117127 149931 117161 149959
rect 117189 149931 117224 149959
rect 117064 149897 117224 149931
rect 117064 149869 117099 149897
rect 117127 149869 117161 149897
rect 117189 149869 117224 149897
rect 117064 149835 117224 149869
rect 117064 149807 117099 149835
rect 117127 149807 117161 149835
rect 117189 149807 117224 149835
rect 117064 149773 117224 149807
rect 117064 149745 117099 149773
rect 117127 149745 117161 149773
rect 117189 149745 117224 149773
rect 117064 149728 117224 149745
rect 132424 149959 132584 149976
rect 132424 149931 132459 149959
rect 132487 149931 132521 149959
rect 132549 149931 132584 149959
rect 132424 149897 132584 149931
rect 132424 149869 132459 149897
rect 132487 149869 132521 149897
rect 132549 149869 132584 149897
rect 132424 149835 132584 149869
rect 132424 149807 132459 149835
rect 132487 149807 132521 149835
rect 132549 149807 132584 149835
rect 132424 149773 132584 149807
rect 132424 149745 132459 149773
rect 132487 149745 132521 149773
rect 132549 149745 132584 149773
rect 132424 149728 132584 149745
rect 147784 149959 147944 149976
rect 147784 149931 147819 149959
rect 147847 149931 147881 149959
rect 147909 149931 147944 149959
rect 147784 149897 147944 149931
rect 147784 149869 147819 149897
rect 147847 149869 147881 149897
rect 147909 149869 147944 149897
rect 147784 149835 147944 149869
rect 147784 149807 147819 149835
rect 147847 149807 147881 149835
rect 147909 149807 147944 149835
rect 147784 149773 147944 149807
rect 147784 149745 147819 149773
rect 147847 149745 147881 149773
rect 147909 149745 147944 149773
rect 147784 149728 147944 149745
rect 163144 149959 163304 149976
rect 163144 149931 163179 149959
rect 163207 149931 163241 149959
rect 163269 149931 163304 149959
rect 163144 149897 163304 149931
rect 163144 149869 163179 149897
rect 163207 149869 163241 149897
rect 163269 149869 163304 149897
rect 163144 149835 163304 149869
rect 163144 149807 163179 149835
rect 163207 149807 163241 149835
rect 163269 149807 163304 149835
rect 163144 149773 163304 149807
rect 163144 149745 163179 149773
rect 163207 149745 163241 149773
rect 163269 149745 163304 149773
rect 163144 149728 163304 149745
rect 178504 149959 178664 149976
rect 178504 149931 178539 149959
rect 178567 149931 178601 149959
rect 178629 149931 178664 149959
rect 178504 149897 178664 149931
rect 178504 149869 178539 149897
rect 178567 149869 178601 149897
rect 178629 149869 178664 149897
rect 178504 149835 178664 149869
rect 178504 149807 178539 149835
rect 178567 149807 178601 149835
rect 178629 149807 178664 149835
rect 178504 149773 178664 149807
rect 178504 149745 178539 149773
rect 178567 149745 178601 149773
rect 178629 149745 178664 149773
rect 178504 149728 178664 149745
rect 193864 149959 194024 149976
rect 193864 149931 193899 149959
rect 193927 149931 193961 149959
rect 193989 149931 194024 149959
rect 193864 149897 194024 149931
rect 193864 149869 193899 149897
rect 193927 149869 193961 149897
rect 193989 149869 194024 149897
rect 193864 149835 194024 149869
rect 193864 149807 193899 149835
rect 193927 149807 193961 149835
rect 193989 149807 194024 149835
rect 193864 149773 194024 149807
rect 193864 149745 193899 149773
rect 193927 149745 193961 149773
rect 193989 149745 194024 149773
rect 193864 149728 194024 149745
rect 209224 149959 209384 149976
rect 209224 149931 209259 149959
rect 209287 149931 209321 149959
rect 209349 149931 209384 149959
rect 209224 149897 209384 149931
rect 209224 149869 209259 149897
rect 209287 149869 209321 149897
rect 209349 149869 209384 149897
rect 209224 149835 209384 149869
rect 209224 149807 209259 149835
rect 209287 149807 209321 149835
rect 209349 149807 209384 149835
rect 209224 149773 209384 149807
rect 209224 149745 209259 149773
rect 209287 149745 209321 149773
rect 209349 149745 209384 149773
rect 209224 149728 209384 149745
rect 224584 149959 224744 149976
rect 224584 149931 224619 149959
rect 224647 149931 224681 149959
rect 224709 149931 224744 149959
rect 224584 149897 224744 149931
rect 224584 149869 224619 149897
rect 224647 149869 224681 149897
rect 224709 149869 224744 149897
rect 224584 149835 224744 149869
rect 224584 149807 224619 149835
rect 224647 149807 224681 149835
rect 224709 149807 224744 149835
rect 224584 149773 224744 149807
rect 224584 149745 224619 149773
rect 224647 149745 224681 149773
rect 224709 149745 224744 149773
rect 224584 149728 224744 149745
rect 239944 149959 240104 149976
rect 239944 149931 239979 149959
rect 240007 149931 240041 149959
rect 240069 149931 240104 149959
rect 239944 149897 240104 149931
rect 239944 149869 239979 149897
rect 240007 149869 240041 149897
rect 240069 149869 240104 149897
rect 239944 149835 240104 149869
rect 239944 149807 239979 149835
rect 240007 149807 240041 149835
rect 240069 149807 240104 149835
rect 239944 149773 240104 149807
rect 239944 149745 239979 149773
rect 240007 149745 240041 149773
rect 240069 149745 240104 149773
rect 239944 149728 240104 149745
rect 32584 146959 32744 146976
rect 32584 146931 32619 146959
rect 32647 146931 32681 146959
rect 32709 146931 32744 146959
rect 32584 146897 32744 146931
rect 32584 146869 32619 146897
rect 32647 146869 32681 146897
rect 32709 146869 32744 146897
rect 32584 146835 32744 146869
rect 32584 146807 32619 146835
rect 32647 146807 32681 146835
rect 32709 146807 32744 146835
rect 32584 146773 32744 146807
rect 32584 146745 32619 146773
rect 32647 146745 32681 146773
rect 32709 146745 32744 146773
rect 32584 146728 32744 146745
rect 47944 146959 48104 146976
rect 47944 146931 47979 146959
rect 48007 146931 48041 146959
rect 48069 146931 48104 146959
rect 47944 146897 48104 146931
rect 47944 146869 47979 146897
rect 48007 146869 48041 146897
rect 48069 146869 48104 146897
rect 47944 146835 48104 146869
rect 47944 146807 47979 146835
rect 48007 146807 48041 146835
rect 48069 146807 48104 146835
rect 47944 146773 48104 146807
rect 47944 146745 47979 146773
rect 48007 146745 48041 146773
rect 48069 146745 48104 146773
rect 47944 146728 48104 146745
rect 63304 146959 63464 146976
rect 63304 146931 63339 146959
rect 63367 146931 63401 146959
rect 63429 146931 63464 146959
rect 63304 146897 63464 146931
rect 63304 146869 63339 146897
rect 63367 146869 63401 146897
rect 63429 146869 63464 146897
rect 63304 146835 63464 146869
rect 63304 146807 63339 146835
rect 63367 146807 63401 146835
rect 63429 146807 63464 146835
rect 63304 146773 63464 146807
rect 63304 146745 63339 146773
rect 63367 146745 63401 146773
rect 63429 146745 63464 146773
rect 63304 146728 63464 146745
rect 78664 146959 78824 146976
rect 78664 146931 78699 146959
rect 78727 146931 78761 146959
rect 78789 146931 78824 146959
rect 78664 146897 78824 146931
rect 78664 146869 78699 146897
rect 78727 146869 78761 146897
rect 78789 146869 78824 146897
rect 78664 146835 78824 146869
rect 78664 146807 78699 146835
rect 78727 146807 78761 146835
rect 78789 146807 78824 146835
rect 78664 146773 78824 146807
rect 78664 146745 78699 146773
rect 78727 146745 78761 146773
rect 78789 146745 78824 146773
rect 78664 146728 78824 146745
rect 94024 146959 94184 146976
rect 94024 146931 94059 146959
rect 94087 146931 94121 146959
rect 94149 146931 94184 146959
rect 94024 146897 94184 146931
rect 94024 146869 94059 146897
rect 94087 146869 94121 146897
rect 94149 146869 94184 146897
rect 94024 146835 94184 146869
rect 94024 146807 94059 146835
rect 94087 146807 94121 146835
rect 94149 146807 94184 146835
rect 94024 146773 94184 146807
rect 94024 146745 94059 146773
rect 94087 146745 94121 146773
rect 94149 146745 94184 146773
rect 94024 146728 94184 146745
rect 109384 146959 109544 146976
rect 109384 146931 109419 146959
rect 109447 146931 109481 146959
rect 109509 146931 109544 146959
rect 109384 146897 109544 146931
rect 109384 146869 109419 146897
rect 109447 146869 109481 146897
rect 109509 146869 109544 146897
rect 109384 146835 109544 146869
rect 109384 146807 109419 146835
rect 109447 146807 109481 146835
rect 109509 146807 109544 146835
rect 109384 146773 109544 146807
rect 109384 146745 109419 146773
rect 109447 146745 109481 146773
rect 109509 146745 109544 146773
rect 109384 146728 109544 146745
rect 124744 146959 124904 146976
rect 124744 146931 124779 146959
rect 124807 146931 124841 146959
rect 124869 146931 124904 146959
rect 124744 146897 124904 146931
rect 124744 146869 124779 146897
rect 124807 146869 124841 146897
rect 124869 146869 124904 146897
rect 124744 146835 124904 146869
rect 124744 146807 124779 146835
rect 124807 146807 124841 146835
rect 124869 146807 124904 146835
rect 124744 146773 124904 146807
rect 124744 146745 124779 146773
rect 124807 146745 124841 146773
rect 124869 146745 124904 146773
rect 124744 146728 124904 146745
rect 140104 146959 140264 146976
rect 140104 146931 140139 146959
rect 140167 146931 140201 146959
rect 140229 146931 140264 146959
rect 140104 146897 140264 146931
rect 140104 146869 140139 146897
rect 140167 146869 140201 146897
rect 140229 146869 140264 146897
rect 140104 146835 140264 146869
rect 140104 146807 140139 146835
rect 140167 146807 140201 146835
rect 140229 146807 140264 146835
rect 140104 146773 140264 146807
rect 140104 146745 140139 146773
rect 140167 146745 140201 146773
rect 140229 146745 140264 146773
rect 140104 146728 140264 146745
rect 155464 146959 155624 146976
rect 155464 146931 155499 146959
rect 155527 146931 155561 146959
rect 155589 146931 155624 146959
rect 155464 146897 155624 146931
rect 155464 146869 155499 146897
rect 155527 146869 155561 146897
rect 155589 146869 155624 146897
rect 155464 146835 155624 146869
rect 155464 146807 155499 146835
rect 155527 146807 155561 146835
rect 155589 146807 155624 146835
rect 155464 146773 155624 146807
rect 155464 146745 155499 146773
rect 155527 146745 155561 146773
rect 155589 146745 155624 146773
rect 155464 146728 155624 146745
rect 170824 146959 170984 146976
rect 170824 146931 170859 146959
rect 170887 146931 170921 146959
rect 170949 146931 170984 146959
rect 170824 146897 170984 146931
rect 170824 146869 170859 146897
rect 170887 146869 170921 146897
rect 170949 146869 170984 146897
rect 170824 146835 170984 146869
rect 170824 146807 170859 146835
rect 170887 146807 170921 146835
rect 170949 146807 170984 146835
rect 170824 146773 170984 146807
rect 170824 146745 170859 146773
rect 170887 146745 170921 146773
rect 170949 146745 170984 146773
rect 170824 146728 170984 146745
rect 186184 146959 186344 146976
rect 186184 146931 186219 146959
rect 186247 146931 186281 146959
rect 186309 146931 186344 146959
rect 186184 146897 186344 146931
rect 186184 146869 186219 146897
rect 186247 146869 186281 146897
rect 186309 146869 186344 146897
rect 186184 146835 186344 146869
rect 186184 146807 186219 146835
rect 186247 146807 186281 146835
rect 186309 146807 186344 146835
rect 186184 146773 186344 146807
rect 186184 146745 186219 146773
rect 186247 146745 186281 146773
rect 186309 146745 186344 146773
rect 186184 146728 186344 146745
rect 201544 146959 201704 146976
rect 201544 146931 201579 146959
rect 201607 146931 201641 146959
rect 201669 146931 201704 146959
rect 201544 146897 201704 146931
rect 201544 146869 201579 146897
rect 201607 146869 201641 146897
rect 201669 146869 201704 146897
rect 201544 146835 201704 146869
rect 201544 146807 201579 146835
rect 201607 146807 201641 146835
rect 201669 146807 201704 146835
rect 201544 146773 201704 146807
rect 201544 146745 201579 146773
rect 201607 146745 201641 146773
rect 201669 146745 201704 146773
rect 201544 146728 201704 146745
rect 216904 146959 217064 146976
rect 216904 146931 216939 146959
rect 216967 146931 217001 146959
rect 217029 146931 217064 146959
rect 216904 146897 217064 146931
rect 216904 146869 216939 146897
rect 216967 146869 217001 146897
rect 217029 146869 217064 146897
rect 216904 146835 217064 146869
rect 216904 146807 216939 146835
rect 216967 146807 217001 146835
rect 217029 146807 217064 146835
rect 216904 146773 217064 146807
rect 216904 146745 216939 146773
rect 216967 146745 217001 146773
rect 217029 146745 217064 146773
rect 216904 146728 217064 146745
rect 232264 146959 232424 146976
rect 232264 146931 232299 146959
rect 232327 146931 232361 146959
rect 232389 146931 232424 146959
rect 232264 146897 232424 146931
rect 232264 146869 232299 146897
rect 232327 146869 232361 146897
rect 232389 146869 232424 146897
rect 232264 146835 232424 146869
rect 232264 146807 232299 146835
rect 232327 146807 232361 146835
rect 232389 146807 232424 146835
rect 232264 146773 232424 146807
rect 232264 146745 232299 146773
rect 232327 146745 232361 146773
rect 232389 146745 232424 146773
rect 232264 146728 232424 146745
rect 247624 146959 247784 146976
rect 247624 146931 247659 146959
rect 247687 146931 247721 146959
rect 247749 146931 247784 146959
rect 247624 146897 247784 146931
rect 247624 146869 247659 146897
rect 247687 146869 247721 146897
rect 247749 146869 247784 146897
rect 247624 146835 247784 146869
rect 247624 146807 247659 146835
rect 247687 146807 247721 146835
rect 247749 146807 247784 146835
rect 247624 146773 247784 146807
rect 247624 146745 247659 146773
rect 247687 146745 247721 146773
rect 247749 146745 247784 146773
rect 247624 146728 247784 146745
rect 254529 146959 254839 155745
rect 254529 146931 254577 146959
rect 254605 146931 254639 146959
rect 254667 146931 254701 146959
rect 254729 146931 254763 146959
rect 254791 146931 254839 146959
rect 254529 146897 254839 146931
rect 254529 146869 254577 146897
rect 254605 146869 254639 146897
rect 254667 146869 254701 146897
rect 254729 146869 254763 146897
rect 254791 146869 254839 146897
rect 254529 146835 254839 146869
rect 254529 146807 254577 146835
rect 254605 146807 254639 146835
rect 254667 146807 254701 146835
rect 254729 146807 254763 146835
rect 254791 146807 254839 146835
rect 254529 146773 254839 146807
rect 254529 146745 254577 146773
rect 254605 146745 254639 146773
rect 254667 146745 254701 146773
rect 254729 146745 254763 146773
rect 254791 146745 254839 146773
rect 31389 140931 31437 140959
rect 31465 140931 31499 140959
rect 31527 140931 31561 140959
rect 31589 140931 31623 140959
rect 31651 140931 31699 140959
rect 31389 140897 31699 140931
rect 31389 140869 31437 140897
rect 31465 140869 31499 140897
rect 31527 140869 31561 140897
rect 31589 140869 31623 140897
rect 31651 140869 31699 140897
rect 31389 140835 31699 140869
rect 31389 140807 31437 140835
rect 31465 140807 31499 140835
rect 31527 140807 31561 140835
rect 31589 140807 31623 140835
rect 31651 140807 31699 140835
rect 31389 140773 31699 140807
rect 31389 140745 31437 140773
rect 31465 140745 31499 140773
rect 31527 140745 31561 140773
rect 31589 140745 31623 140773
rect 31651 140745 31699 140773
rect 31389 131959 31699 140745
rect 40264 140959 40424 140976
rect 40264 140931 40299 140959
rect 40327 140931 40361 140959
rect 40389 140931 40424 140959
rect 40264 140897 40424 140931
rect 40264 140869 40299 140897
rect 40327 140869 40361 140897
rect 40389 140869 40424 140897
rect 40264 140835 40424 140869
rect 40264 140807 40299 140835
rect 40327 140807 40361 140835
rect 40389 140807 40424 140835
rect 40264 140773 40424 140807
rect 40264 140745 40299 140773
rect 40327 140745 40361 140773
rect 40389 140745 40424 140773
rect 40264 140728 40424 140745
rect 55624 140959 55784 140976
rect 55624 140931 55659 140959
rect 55687 140931 55721 140959
rect 55749 140931 55784 140959
rect 55624 140897 55784 140931
rect 55624 140869 55659 140897
rect 55687 140869 55721 140897
rect 55749 140869 55784 140897
rect 55624 140835 55784 140869
rect 55624 140807 55659 140835
rect 55687 140807 55721 140835
rect 55749 140807 55784 140835
rect 55624 140773 55784 140807
rect 55624 140745 55659 140773
rect 55687 140745 55721 140773
rect 55749 140745 55784 140773
rect 55624 140728 55784 140745
rect 70984 140959 71144 140976
rect 70984 140931 71019 140959
rect 71047 140931 71081 140959
rect 71109 140931 71144 140959
rect 70984 140897 71144 140931
rect 70984 140869 71019 140897
rect 71047 140869 71081 140897
rect 71109 140869 71144 140897
rect 70984 140835 71144 140869
rect 70984 140807 71019 140835
rect 71047 140807 71081 140835
rect 71109 140807 71144 140835
rect 70984 140773 71144 140807
rect 70984 140745 71019 140773
rect 71047 140745 71081 140773
rect 71109 140745 71144 140773
rect 70984 140728 71144 140745
rect 86344 140959 86504 140976
rect 86344 140931 86379 140959
rect 86407 140931 86441 140959
rect 86469 140931 86504 140959
rect 86344 140897 86504 140931
rect 86344 140869 86379 140897
rect 86407 140869 86441 140897
rect 86469 140869 86504 140897
rect 86344 140835 86504 140869
rect 86344 140807 86379 140835
rect 86407 140807 86441 140835
rect 86469 140807 86504 140835
rect 86344 140773 86504 140807
rect 86344 140745 86379 140773
rect 86407 140745 86441 140773
rect 86469 140745 86504 140773
rect 86344 140728 86504 140745
rect 101704 140959 101864 140976
rect 101704 140931 101739 140959
rect 101767 140931 101801 140959
rect 101829 140931 101864 140959
rect 101704 140897 101864 140931
rect 101704 140869 101739 140897
rect 101767 140869 101801 140897
rect 101829 140869 101864 140897
rect 101704 140835 101864 140869
rect 101704 140807 101739 140835
rect 101767 140807 101801 140835
rect 101829 140807 101864 140835
rect 101704 140773 101864 140807
rect 101704 140745 101739 140773
rect 101767 140745 101801 140773
rect 101829 140745 101864 140773
rect 101704 140728 101864 140745
rect 117064 140959 117224 140976
rect 117064 140931 117099 140959
rect 117127 140931 117161 140959
rect 117189 140931 117224 140959
rect 117064 140897 117224 140931
rect 117064 140869 117099 140897
rect 117127 140869 117161 140897
rect 117189 140869 117224 140897
rect 117064 140835 117224 140869
rect 117064 140807 117099 140835
rect 117127 140807 117161 140835
rect 117189 140807 117224 140835
rect 117064 140773 117224 140807
rect 117064 140745 117099 140773
rect 117127 140745 117161 140773
rect 117189 140745 117224 140773
rect 117064 140728 117224 140745
rect 132424 140959 132584 140976
rect 132424 140931 132459 140959
rect 132487 140931 132521 140959
rect 132549 140931 132584 140959
rect 132424 140897 132584 140931
rect 132424 140869 132459 140897
rect 132487 140869 132521 140897
rect 132549 140869 132584 140897
rect 132424 140835 132584 140869
rect 132424 140807 132459 140835
rect 132487 140807 132521 140835
rect 132549 140807 132584 140835
rect 132424 140773 132584 140807
rect 132424 140745 132459 140773
rect 132487 140745 132521 140773
rect 132549 140745 132584 140773
rect 132424 140728 132584 140745
rect 147784 140959 147944 140976
rect 147784 140931 147819 140959
rect 147847 140931 147881 140959
rect 147909 140931 147944 140959
rect 147784 140897 147944 140931
rect 147784 140869 147819 140897
rect 147847 140869 147881 140897
rect 147909 140869 147944 140897
rect 147784 140835 147944 140869
rect 147784 140807 147819 140835
rect 147847 140807 147881 140835
rect 147909 140807 147944 140835
rect 147784 140773 147944 140807
rect 147784 140745 147819 140773
rect 147847 140745 147881 140773
rect 147909 140745 147944 140773
rect 147784 140728 147944 140745
rect 163144 140959 163304 140976
rect 163144 140931 163179 140959
rect 163207 140931 163241 140959
rect 163269 140931 163304 140959
rect 163144 140897 163304 140931
rect 163144 140869 163179 140897
rect 163207 140869 163241 140897
rect 163269 140869 163304 140897
rect 163144 140835 163304 140869
rect 163144 140807 163179 140835
rect 163207 140807 163241 140835
rect 163269 140807 163304 140835
rect 163144 140773 163304 140807
rect 163144 140745 163179 140773
rect 163207 140745 163241 140773
rect 163269 140745 163304 140773
rect 163144 140728 163304 140745
rect 178504 140959 178664 140976
rect 178504 140931 178539 140959
rect 178567 140931 178601 140959
rect 178629 140931 178664 140959
rect 178504 140897 178664 140931
rect 178504 140869 178539 140897
rect 178567 140869 178601 140897
rect 178629 140869 178664 140897
rect 178504 140835 178664 140869
rect 178504 140807 178539 140835
rect 178567 140807 178601 140835
rect 178629 140807 178664 140835
rect 178504 140773 178664 140807
rect 178504 140745 178539 140773
rect 178567 140745 178601 140773
rect 178629 140745 178664 140773
rect 178504 140728 178664 140745
rect 193864 140959 194024 140976
rect 193864 140931 193899 140959
rect 193927 140931 193961 140959
rect 193989 140931 194024 140959
rect 193864 140897 194024 140931
rect 193864 140869 193899 140897
rect 193927 140869 193961 140897
rect 193989 140869 194024 140897
rect 193864 140835 194024 140869
rect 193864 140807 193899 140835
rect 193927 140807 193961 140835
rect 193989 140807 194024 140835
rect 193864 140773 194024 140807
rect 193864 140745 193899 140773
rect 193927 140745 193961 140773
rect 193989 140745 194024 140773
rect 193864 140728 194024 140745
rect 209224 140959 209384 140976
rect 209224 140931 209259 140959
rect 209287 140931 209321 140959
rect 209349 140931 209384 140959
rect 209224 140897 209384 140931
rect 209224 140869 209259 140897
rect 209287 140869 209321 140897
rect 209349 140869 209384 140897
rect 209224 140835 209384 140869
rect 209224 140807 209259 140835
rect 209287 140807 209321 140835
rect 209349 140807 209384 140835
rect 209224 140773 209384 140807
rect 209224 140745 209259 140773
rect 209287 140745 209321 140773
rect 209349 140745 209384 140773
rect 209224 140728 209384 140745
rect 224584 140959 224744 140976
rect 224584 140931 224619 140959
rect 224647 140931 224681 140959
rect 224709 140931 224744 140959
rect 224584 140897 224744 140931
rect 224584 140869 224619 140897
rect 224647 140869 224681 140897
rect 224709 140869 224744 140897
rect 224584 140835 224744 140869
rect 224584 140807 224619 140835
rect 224647 140807 224681 140835
rect 224709 140807 224744 140835
rect 224584 140773 224744 140807
rect 224584 140745 224619 140773
rect 224647 140745 224681 140773
rect 224709 140745 224744 140773
rect 224584 140728 224744 140745
rect 239944 140959 240104 140976
rect 239944 140931 239979 140959
rect 240007 140931 240041 140959
rect 240069 140931 240104 140959
rect 239944 140897 240104 140931
rect 239944 140869 239979 140897
rect 240007 140869 240041 140897
rect 240069 140869 240104 140897
rect 239944 140835 240104 140869
rect 239944 140807 239979 140835
rect 240007 140807 240041 140835
rect 240069 140807 240104 140835
rect 239944 140773 240104 140807
rect 239944 140745 239979 140773
rect 240007 140745 240041 140773
rect 240069 140745 240104 140773
rect 239944 140728 240104 140745
rect 32584 137959 32744 137976
rect 32584 137931 32619 137959
rect 32647 137931 32681 137959
rect 32709 137931 32744 137959
rect 32584 137897 32744 137931
rect 32584 137869 32619 137897
rect 32647 137869 32681 137897
rect 32709 137869 32744 137897
rect 32584 137835 32744 137869
rect 32584 137807 32619 137835
rect 32647 137807 32681 137835
rect 32709 137807 32744 137835
rect 32584 137773 32744 137807
rect 32584 137745 32619 137773
rect 32647 137745 32681 137773
rect 32709 137745 32744 137773
rect 32584 137728 32744 137745
rect 47944 137959 48104 137976
rect 47944 137931 47979 137959
rect 48007 137931 48041 137959
rect 48069 137931 48104 137959
rect 47944 137897 48104 137931
rect 47944 137869 47979 137897
rect 48007 137869 48041 137897
rect 48069 137869 48104 137897
rect 47944 137835 48104 137869
rect 47944 137807 47979 137835
rect 48007 137807 48041 137835
rect 48069 137807 48104 137835
rect 47944 137773 48104 137807
rect 47944 137745 47979 137773
rect 48007 137745 48041 137773
rect 48069 137745 48104 137773
rect 47944 137728 48104 137745
rect 63304 137959 63464 137976
rect 63304 137931 63339 137959
rect 63367 137931 63401 137959
rect 63429 137931 63464 137959
rect 63304 137897 63464 137931
rect 63304 137869 63339 137897
rect 63367 137869 63401 137897
rect 63429 137869 63464 137897
rect 63304 137835 63464 137869
rect 63304 137807 63339 137835
rect 63367 137807 63401 137835
rect 63429 137807 63464 137835
rect 63304 137773 63464 137807
rect 63304 137745 63339 137773
rect 63367 137745 63401 137773
rect 63429 137745 63464 137773
rect 63304 137728 63464 137745
rect 78664 137959 78824 137976
rect 78664 137931 78699 137959
rect 78727 137931 78761 137959
rect 78789 137931 78824 137959
rect 78664 137897 78824 137931
rect 78664 137869 78699 137897
rect 78727 137869 78761 137897
rect 78789 137869 78824 137897
rect 78664 137835 78824 137869
rect 78664 137807 78699 137835
rect 78727 137807 78761 137835
rect 78789 137807 78824 137835
rect 78664 137773 78824 137807
rect 78664 137745 78699 137773
rect 78727 137745 78761 137773
rect 78789 137745 78824 137773
rect 78664 137728 78824 137745
rect 94024 137959 94184 137976
rect 94024 137931 94059 137959
rect 94087 137931 94121 137959
rect 94149 137931 94184 137959
rect 94024 137897 94184 137931
rect 94024 137869 94059 137897
rect 94087 137869 94121 137897
rect 94149 137869 94184 137897
rect 94024 137835 94184 137869
rect 94024 137807 94059 137835
rect 94087 137807 94121 137835
rect 94149 137807 94184 137835
rect 94024 137773 94184 137807
rect 94024 137745 94059 137773
rect 94087 137745 94121 137773
rect 94149 137745 94184 137773
rect 94024 137728 94184 137745
rect 109384 137959 109544 137976
rect 109384 137931 109419 137959
rect 109447 137931 109481 137959
rect 109509 137931 109544 137959
rect 109384 137897 109544 137931
rect 109384 137869 109419 137897
rect 109447 137869 109481 137897
rect 109509 137869 109544 137897
rect 109384 137835 109544 137869
rect 109384 137807 109419 137835
rect 109447 137807 109481 137835
rect 109509 137807 109544 137835
rect 109384 137773 109544 137807
rect 109384 137745 109419 137773
rect 109447 137745 109481 137773
rect 109509 137745 109544 137773
rect 109384 137728 109544 137745
rect 124744 137959 124904 137976
rect 124744 137931 124779 137959
rect 124807 137931 124841 137959
rect 124869 137931 124904 137959
rect 124744 137897 124904 137931
rect 124744 137869 124779 137897
rect 124807 137869 124841 137897
rect 124869 137869 124904 137897
rect 124744 137835 124904 137869
rect 124744 137807 124779 137835
rect 124807 137807 124841 137835
rect 124869 137807 124904 137835
rect 124744 137773 124904 137807
rect 124744 137745 124779 137773
rect 124807 137745 124841 137773
rect 124869 137745 124904 137773
rect 124744 137728 124904 137745
rect 140104 137959 140264 137976
rect 140104 137931 140139 137959
rect 140167 137931 140201 137959
rect 140229 137931 140264 137959
rect 140104 137897 140264 137931
rect 140104 137869 140139 137897
rect 140167 137869 140201 137897
rect 140229 137869 140264 137897
rect 140104 137835 140264 137869
rect 140104 137807 140139 137835
rect 140167 137807 140201 137835
rect 140229 137807 140264 137835
rect 140104 137773 140264 137807
rect 140104 137745 140139 137773
rect 140167 137745 140201 137773
rect 140229 137745 140264 137773
rect 140104 137728 140264 137745
rect 155464 137959 155624 137976
rect 155464 137931 155499 137959
rect 155527 137931 155561 137959
rect 155589 137931 155624 137959
rect 155464 137897 155624 137931
rect 155464 137869 155499 137897
rect 155527 137869 155561 137897
rect 155589 137869 155624 137897
rect 155464 137835 155624 137869
rect 155464 137807 155499 137835
rect 155527 137807 155561 137835
rect 155589 137807 155624 137835
rect 155464 137773 155624 137807
rect 155464 137745 155499 137773
rect 155527 137745 155561 137773
rect 155589 137745 155624 137773
rect 155464 137728 155624 137745
rect 170824 137959 170984 137976
rect 170824 137931 170859 137959
rect 170887 137931 170921 137959
rect 170949 137931 170984 137959
rect 170824 137897 170984 137931
rect 170824 137869 170859 137897
rect 170887 137869 170921 137897
rect 170949 137869 170984 137897
rect 170824 137835 170984 137869
rect 170824 137807 170859 137835
rect 170887 137807 170921 137835
rect 170949 137807 170984 137835
rect 170824 137773 170984 137807
rect 170824 137745 170859 137773
rect 170887 137745 170921 137773
rect 170949 137745 170984 137773
rect 170824 137728 170984 137745
rect 186184 137959 186344 137976
rect 186184 137931 186219 137959
rect 186247 137931 186281 137959
rect 186309 137931 186344 137959
rect 186184 137897 186344 137931
rect 186184 137869 186219 137897
rect 186247 137869 186281 137897
rect 186309 137869 186344 137897
rect 186184 137835 186344 137869
rect 186184 137807 186219 137835
rect 186247 137807 186281 137835
rect 186309 137807 186344 137835
rect 186184 137773 186344 137807
rect 186184 137745 186219 137773
rect 186247 137745 186281 137773
rect 186309 137745 186344 137773
rect 186184 137728 186344 137745
rect 201544 137959 201704 137976
rect 201544 137931 201579 137959
rect 201607 137931 201641 137959
rect 201669 137931 201704 137959
rect 201544 137897 201704 137931
rect 201544 137869 201579 137897
rect 201607 137869 201641 137897
rect 201669 137869 201704 137897
rect 201544 137835 201704 137869
rect 201544 137807 201579 137835
rect 201607 137807 201641 137835
rect 201669 137807 201704 137835
rect 201544 137773 201704 137807
rect 201544 137745 201579 137773
rect 201607 137745 201641 137773
rect 201669 137745 201704 137773
rect 201544 137728 201704 137745
rect 216904 137959 217064 137976
rect 216904 137931 216939 137959
rect 216967 137931 217001 137959
rect 217029 137931 217064 137959
rect 216904 137897 217064 137931
rect 216904 137869 216939 137897
rect 216967 137869 217001 137897
rect 217029 137869 217064 137897
rect 216904 137835 217064 137869
rect 216904 137807 216939 137835
rect 216967 137807 217001 137835
rect 217029 137807 217064 137835
rect 216904 137773 217064 137807
rect 216904 137745 216939 137773
rect 216967 137745 217001 137773
rect 217029 137745 217064 137773
rect 216904 137728 217064 137745
rect 232264 137959 232424 137976
rect 232264 137931 232299 137959
rect 232327 137931 232361 137959
rect 232389 137931 232424 137959
rect 232264 137897 232424 137931
rect 232264 137869 232299 137897
rect 232327 137869 232361 137897
rect 232389 137869 232424 137897
rect 232264 137835 232424 137869
rect 232264 137807 232299 137835
rect 232327 137807 232361 137835
rect 232389 137807 232424 137835
rect 232264 137773 232424 137807
rect 232264 137745 232299 137773
rect 232327 137745 232361 137773
rect 232389 137745 232424 137773
rect 232264 137728 232424 137745
rect 247624 137959 247784 137976
rect 247624 137931 247659 137959
rect 247687 137931 247721 137959
rect 247749 137931 247784 137959
rect 247624 137897 247784 137931
rect 247624 137869 247659 137897
rect 247687 137869 247721 137897
rect 247749 137869 247784 137897
rect 247624 137835 247784 137869
rect 247624 137807 247659 137835
rect 247687 137807 247721 137835
rect 247749 137807 247784 137835
rect 247624 137773 247784 137807
rect 247624 137745 247659 137773
rect 247687 137745 247721 137773
rect 247749 137745 247784 137773
rect 247624 137728 247784 137745
rect 254529 137959 254839 146745
rect 254529 137931 254577 137959
rect 254605 137931 254639 137959
rect 254667 137931 254701 137959
rect 254729 137931 254763 137959
rect 254791 137931 254839 137959
rect 254529 137897 254839 137931
rect 254529 137869 254577 137897
rect 254605 137869 254639 137897
rect 254667 137869 254701 137897
rect 254729 137869 254763 137897
rect 254791 137869 254839 137897
rect 254529 137835 254839 137869
rect 254529 137807 254577 137835
rect 254605 137807 254639 137835
rect 254667 137807 254701 137835
rect 254729 137807 254763 137835
rect 254791 137807 254839 137835
rect 254529 137773 254839 137807
rect 254529 137745 254577 137773
rect 254605 137745 254639 137773
rect 254667 137745 254701 137773
rect 254729 137745 254763 137773
rect 254791 137745 254839 137773
rect 31389 131931 31437 131959
rect 31465 131931 31499 131959
rect 31527 131931 31561 131959
rect 31589 131931 31623 131959
rect 31651 131931 31699 131959
rect 31389 131897 31699 131931
rect 31389 131869 31437 131897
rect 31465 131869 31499 131897
rect 31527 131869 31561 131897
rect 31589 131869 31623 131897
rect 31651 131869 31699 131897
rect 31389 131835 31699 131869
rect 31389 131807 31437 131835
rect 31465 131807 31499 131835
rect 31527 131807 31561 131835
rect 31589 131807 31623 131835
rect 31651 131807 31699 131835
rect 31389 131773 31699 131807
rect 31389 131745 31437 131773
rect 31465 131745 31499 131773
rect 31527 131745 31561 131773
rect 31589 131745 31623 131773
rect 31651 131745 31699 131773
rect 31389 122959 31699 131745
rect 40264 131959 40424 131976
rect 40264 131931 40299 131959
rect 40327 131931 40361 131959
rect 40389 131931 40424 131959
rect 40264 131897 40424 131931
rect 40264 131869 40299 131897
rect 40327 131869 40361 131897
rect 40389 131869 40424 131897
rect 40264 131835 40424 131869
rect 40264 131807 40299 131835
rect 40327 131807 40361 131835
rect 40389 131807 40424 131835
rect 40264 131773 40424 131807
rect 40264 131745 40299 131773
rect 40327 131745 40361 131773
rect 40389 131745 40424 131773
rect 40264 131728 40424 131745
rect 55624 131959 55784 131976
rect 55624 131931 55659 131959
rect 55687 131931 55721 131959
rect 55749 131931 55784 131959
rect 55624 131897 55784 131931
rect 55624 131869 55659 131897
rect 55687 131869 55721 131897
rect 55749 131869 55784 131897
rect 55624 131835 55784 131869
rect 55624 131807 55659 131835
rect 55687 131807 55721 131835
rect 55749 131807 55784 131835
rect 55624 131773 55784 131807
rect 55624 131745 55659 131773
rect 55687 131745 55721 131773
rect 55749 131745 55784 131773
rect 55624 131728 55784 131745
rect 70984 131959 71144 131976
rect 70984 131931 71019 131959
rect 71047 131931 71081 131959
rect 71109 131931 71144 131959
rect 70984 131897 71144 131931
rect 70984 131869 71019 131897
rect 71047 131869 71081 131897
rect 71109 131869 71144 131897
rect 70984 131835 71144 131869
rect 70984 131807 71019 131835
rect 71047 131807 71081 131835
rect 71109 131807 71144 131835
rect 70984 131773 71144 131807
rect 70984 131745 71019 131773
rect 71047 131745 71081 131773
rect 71109 131745 71144 131773
rect 70984 131728 71144 131745
rect 86344 131959 86504 131976
rect 86344 131931 86379 131959
rect 86407 131931 86441 131959
rect 86469 131931 86504 131959
rect 86344 131897 86504 131931
rect 86344 131869 86379 131897
rect 86407 131869 86441 131897
rect 86469 131869 86504 131897
rect 86344 131835 86504 131869
rect 86344 131807 86379 131835
rect 86407 131807 86441 131835
rect 86469 131807 86504 131835
rect 86344 131773 86504 131807
rect 86344 131745 86379 131773
rect 86407 131745 86441 131773
rect 86469 131745 86504 131773
rect 86344 131728 86504 131745
rect 101704 131959 101864 131976
rect 101704 131931 101739 131959
rect 101767 131931 101801 131959
rect 101829 131931 101864 131959
rect 101704 131897 101864 131931
rect 101704 131869 101739 131897
rect 101767 131869 101801 131897
rect 101829 131869 101864 131897
rect 101704 131835 101864 131869
rect 101704 131807 101739 131835
rect 101767 131807 101801 131835
rect 101829 131807 101864 131835
rect 101704 131773 101864 131807
rect 101704 131745 101739 131773
rect 101767 131745 101801 131773
rect 101829 131745 101864 131773
rect 101704 131728 101864 131745
rect 117064 131959 117224 131976
rect 117064 131931 117099 131959
rect 117127 131931 117161 131959
rect 117189 131931 117224 131959
rect 117064 131897 117224 131931
rect 117064 131869 117099 131897
rect 117127 131869 117161 131897
rect 117189 131869 117224 131897
rect 117064 131835 117224 131869
rect 117064 131807 117099 131835
rect 117127 131807 117161 131835
rect 117189 131807 117224 131835
rect 117064 131773 117224 131807
rect 117064 131745 117099 131773
rect 117127 131745 117161 131773
rect 117189 131745 117224 131773
rect 117064 131728 117224 131745
rect 132424 131959 132584 131976
rect 132424 131931 132459 131959
rect 132487 131931 132521 131959
rect 132549 131931 132584 131959
rect 132424 131897 132584 131931
rect 132424 131869 132459 131897
rect 132487 131869 132521 131897
rect 132549 131869 132584 131897
rect 132424 131835 132584 131869
rect 132424 131807 132459 131835
rect 132487 131807 132521 131835
rect 132549 131807 132584 131835
rect 132424 131773 132584 131807
rect 132424 131745 132459 131773
rect 132487 131745 132521 131773
rect 132549 131745 132584 131773
rect 132424 131728 132584 131745
rect 147784 131959 147944 131976
rect 147784 131931 147819 131959
rect 147847 131931 147881 131959
rect 147909 131931 147944 131959
rect 147784 131897 147944 131931
rect 147784 131869 147819 131897
rect 147847 131869 147881 131897
rect 147909 131869 147944 131897
rect 147784 131835 147944 131869
rect 147784 131807 147819 131835
rect 147847 131807 147881 131835
rect 147909 131807 147944 131835
rect 147784 131773 147944 131807
rect 147784 131745 147819 131773
rect 147847 131745 147881 131773
rect 147909 131745 147944 131773
rect 147784 131728 147944 131745
rect 163144 131959 163304 131976
rect 163144 131931 163179 131959
rect 163207 131931 163241 131959
rect 163269 131931 163304 131959
rect 163144 131897 163304 131931
rect 163144 131869 163179 131897
rect 163207 131869 163241 131897
rect 163269 131869 163304 131897
rect 163144 131835 163304 131869
rect 163144 131807 163179 131835
rect 163207 131807 163241 131835
rect 163269 131807 163304 131835
rect 163144 131773 163304 131807
rect 163144 131745 163179 131773
rect 163207 131745 163241 131773
rect 163269 131745 163304 131773
rect 163144 131728 163304 131745
rect 178504 131959 178664 131976
rect 178504 131931 178539 131959
rect 178567 131931 178601 131959
rect 178629 131931 178664 131959
rect 178504 131897 178664 131931
rect 178504 131869 178539 131897
rect 178567 131869 178601 131897
rect 178629 131869 178664 131897
rect 178504 131835 178664 131869
rect 178504 131807 178539 131835
rect 178567 131807 178601 131835
rect 178629 131807 178664 131835
rect 178504 131773 178664 131807
rect 178504 131745 178539 131773
rect 178567 131745 178601 131773
rect 178629 131745 178664 131773
rect 178504 131728 178664 131745
rect 193864 131959 194024 131976
rect 193864 131931 193899 131959
rect 193927 131931 193961 131959
rect 193989 131931 194024 131959
rect 193864 131897 194024 131931
rect 193864 131869 193899 131897
rect 193927 131869 193961 131897
rect 193989 131869 194024 131897
rect 193864 131835 194024 131869
rect 193864 131807 193899 131835
rect 193927 131807 193961 131835
rect 193989 131807 194024 131835
rect 193864 131773 194024 131807
rect 193864 131745 193899 131773
rect 193927 131745 193961 131773
rect 193989 131745 194024 131773
rect 193864 131728 194024 131745
rect 209224 131959 209384 131976
rect 209224 131931 209259 131959
rect 209287 131931 209321 131959
rect 209349 131931 209384 131959
rect 209224 131897 209384 131931
rect 209224 131869 209259 131897
rect 209287 131869 209321 131897
rect 209349 131869 209384 131897
rect 209224 131835 209384 131869
rect 209224 131807 209259 131835
rect 209287 131807 209321 131835
rect 209349 131807 209384 131835
rect 209224 131773 209384 131807
rect 209224 131745 209259 131773
rect 209287 131745 209321 131773
rect 209349 131745 209384 131773
rect 209224 131728 209384 131745
rect 224584 131959 224744 131976
rect 224584 131931 224619 131959
rect 224647 131931 224681 131959
rect 224709 131931 224744 131959
rect 224584 131897 224744 131931
rect 224584 131869 224619 131897
rect 224647 131869 224681 131897
rect 224709 131869 224744 131897
rect 224584 131835 224744 131869
rect 224584 131807 224619 131835
rect 224647 131807 224681 131835
rect 224709 131807 224744 131835
rect 224584 131773 224744 131807
rect 224584 131745 224619 131773
rect 224647 131745 224681 131773
rect 224709 131745 224744 131773
rect 224584 131728 224744 131745
rect 239944 131959 240104 131976
rect 239944 131931 239979 131959
rect 240007 131931 240041 131959
rect 240069 131931 240104 131959
rect 239944 131897 240104 131931
rect 239944 131869 239979 131897
rect 240007 131869 240041 131897
rect 240069 131869 240104 131897
rect 239944 131835 240104 131869
rect 239944 131807 239979 131835
rect 240007 131807 240041 131835
rect 240069 131807 240104 131835
rect 239944 131773 240104 131807
rect 239944 131745 239979 131773
rect 240007 131745 240041 131773
rect 240069 131745 240104 131773
rect 239944 131728 240104 131745
rect 32584 128959 32744 128976
rect 32584 128931 32619 128959
rect 32647 128931 32681 128959
rect 32709 128931 32744 128959
rect 32584 128897 32744 128931
rect 32584 128869 32619 128897
rect 32647 128869 32681 128897
rect 32709 128869 32744 128897
rect 32584 128835 32744 128869
rect 32584 128807 32619 128835
rect 32647 128807 32681 128835
rect 32709 128807 32744 128835
rect 32584 128773 32744 128807
rect 32584 128745 32619 128773
rect 32647 128745 32681 128773
rect 32709 128745 32744 128773
rect 32584 128728 32744 128745
rect 47944 128959 48104 128976
rect 47944 128931 47979 128959
rect 48007 128931 48041 128959
rect 48069 128931 48104 128959
rect 47944 128897 48104 128931
rect 47944 128869 47979 128897
rect 48007 128869 48041 128897
rect 48069 128869 48104 128897
rect 47944 128835 48104 128869
rect 47944 128807 47979 128835
rect 48007 128807 48041 128835
rect 48069 128807 48104 128835
rect 47944 128773 48104 128807
rect 47944 128745 47979 128773
rect 48007 128745 48041 128773
rect 48069 128745 48104 128773
rect 47944 128728 48104 128745
rect 63304 128959 63464 128976
rect 63304 128931 63339 128959
rect 63367 128931 63401 128959
rect 63429 128931 63464 128959
rect 63304 128897 63464 128931
rect 63304 128869 63339 128897
rect 63367 128869 63401 128897
rect 63429 128869 63464 128897
rect 63304 128835 63464 128869
rect 63304 128807 63339 128835
rect 63367 128807 63401 128835
rect 63429 128807 63464 128835
rect 63304 128773 63464 128807
rect 63304 128745 63339 128773
rect 63367 128745 63401 128773
rect 63429 128745 63464 128773
rect 63304 128728 63464 128745
rect 78664 128959 78824 128976
rect 78664 128931 78699 128959
rect 78727 128931 78761 128959
rect 78789 128931 78824 128959
rect 78664 128897 78824 128931
rect 78664 128869 78699 128897
rect 78727 128869 78761 128897
rect 78789 128869 78824 128897
rect 78664 128835 78824 128869
rect 78664 128807 78699 128835
rect 78727 128807 78761 128835
rect 78789 128807 78824 128835
rect 78664 128773 78824 128807
rect 78664 128745 78699 128773
rect 78727 128745 78761 128773
rect 78789 128745 78824 128773
rect 78664 128728 78824 128745
rect 94024 128959 94184 128976
rect 94024 128931 94059 128959
rect 94087 128931 94121 128959
rect 94149 128931 94184 128959
rect 94024 128897 94184 128931
rect 94024 128869 94059 128897
rect 94087 128869 94121 128897
rect 94149 128869 94184 128897
rect 94024 128835 94184 128869
rect 94024 128807 94059 128835
rect 94087 128807 94121 128835
rect 94149 128807 94184 128835
rect 94024 128773 94184 128807
rect 94024 128745 94059 128773
rect 94087 128745 94121 128773
rect 94149 128745 94184 128773
rect 94024 128728 94184 128745
rect 109384 128959 109544 128976
rect 109384 128931 109419 128959
rect 109447 128931 109481 128959
rect 109509 128931 109544 128959
rect 109384 128897 109544 128931
rect 109384 128869 109419 128897
rect 109447 128869 109481 128897
rect 109509 128869 109544 128897
rect 109384 128835 109544 128869
rect 109384 128807 109419 128835
rect 109447 128807 109481 128835
rect 109509 128807 109544 128835
rect 109384 128773 109544 128807
rect 109384 128745 109419 128773
rect 109447 128745 109481 128773
rect 109509 128745 109544 128773
rect 109384 128728 109544 128745
rect 124744 128959 124904 128976
rect 124744 128931 124779 128959
rect 124807 128931 124841 128959
rect 124869 128931 124904 128959
rect 124744 128897 124904 128931
rect 124744 128869 124779 128897
rect 124807 128869 124841 128897
rect 124869 128869 124904 128897
rect 124744 128835 124904 128869
rect 124744 128807 124779 128835
rect 124807 128807 124841 128835
rect 124869 128807 124904 128835
rect 124744 128773 124904 128807
rect 124744 128745 124779 128773
rect 124807 128745 124841 128773
rect 124869 128745 124904 128773
rect 124744 128728 124904 128745
rect 140104 128959 140264 128976
rect 140104 128931 140139 128959
rect 140167 128931 140201 128959
rect 140229 128931 140264 128959
rect 140104 128897 140264 128931
rect 140104 128869 140139 128897
rect 140167 128869 140201 128897
rect 140229 128869 140264 128897
rect 140104 128835 140264 128869
rect 140104 128807 140139 128835
rect 140167 128807 140201 128835
rect 140229 128807 140264 128835
rect 140104 128773 140264 128807
rect 140104 128745 140139 128773
rect 140167 128745 140201 128773
rect 140229 128745 140264 128773
rect 140104 128728 140264 128745
rect 155464 128959 155624 128976
rect 155464 128931 155499 128959
rect 155527 128931 155561 128959
rect 155589 128931 155624 128959
rect 155464 128897 155624 128931
rect 155464 128869 155499 128897
rect 155527 128869 155561 128897
rect 155589 128869 155624 128897
rect 155464 128835 155624 128869
rect 155464 128807 155499 128835
rect 155527 128807 155561 128835
rect 155589 128807 155624 128835
rect 155464 128773 155624 128807
rect 155464 128745 155499 128773
rect 155527 128745 155561 128773
rect 155589 128745 155624 128773
rect 155464 128728 155624 128745
rect 170824 128959 170984 128976
rect 170824 128931 170859 128959
rect 170887 128931 170921 128959
rect 170949 128931 170984 128959
rect 170824 128897 170984 128931
rect 170824 128869 170859 128897
rect 170887 128869 170921 128897
rect 170949 128869 170984 128897
rect 170824 128835 170984 128869
rect 170824 128807 170859 128835
rect 170887 128807 170921 128835
rect 170949 128807 170984 128835
rect 170824 128773 170984 128807
rect 170824 128745 170859 128773
rect 170887 128745 170921 128773
rect 170949 128745 170984 128773
rect 170824 128728 170984 128745
rect 186184 128959 186344 128976
rect 186184 128931 186219 128959
rect 186247 128931 186281 128959
rect 186309 128931 186344 128959
rect 186184 128897 186344 128931
rect 186184 128869 186219 128897
rect 186247 128869 186281 128897
rect 186309 128869 186344 128897
rect 186184 128835 186344 128869
rect 186184 128807 186219 128835
rect 186247 128807 186281 128835
rect 186309 128807 186344 128835
rect 186184 128773 186344 128807
rect 186184 128745 186219 128773
rect 186247 128745 186281 128773
rect 186309 128745 186344 128773
rect 186184 128728 186344 128745
rect 201544 128959 201704 128976
rect 201544 128931 201579 128959
rect 201607 128931 201641 128959
rect 201669 128931 201704 128959
rect 201544 128897 201704 128931
rect 201544 128869 201579 128897
rect 201607 128869 201641 128897
rect 201669 128869 201704 128897
rect 201544 128835 201704 128869
rect 201544 128807 201579 128835
rect 201607 128807 201641 128835
rect 201669 128807 201704 128835
rect 201544 128773 201704 128807
rect 201544 128745 201579 128773
rect 201607 128745 201641 128773
rect 201669 128745 201704 128773
rect 201544 128728 201704 128745
rect 216904 128959 217064 128976
rect 216904 128931 216939 128959
rect 216967 128931 217001 128959
rect 217029 128931 217064 128959
rect 216904 128897 217064 128931
rect 216904 128869 216939 128897
rect 216967 128869 217001 128897
rect 217029 128869 217064 128897
rect 216904 128835 217064 128869
rect 216904 128807 216939 128835
rect 216967 128807 217001 128835
rect 217029 128807 217064 128835
rect 216904 128773 217064 128807
rect 216904 128745 216939 128773
rect 216967 128745 217001 128773
rect 217029 128745 217064 128773
rect 216904 128728 217064 128745
rect 232264 128959 232424 128976
rect 232264 128931 232299 128959
rect 232327 128931 232361 128959
rect 232389 128931 232424 128959
rect 232264 128897 232424 128931
rect 232264 128869 232299 128897
rect 232327 128869 232361 128897
rect 232389 128869 232424 128897
rect 232264 128835 232424 128869
rect 232264 128807 232299 128835
rect 232327 128807 232361 128835
rect 232389 128807 232424 128835
rect 232264 128773 232424 128807
rect 232264 128745 232299 128773
rect 232327 128745 232361 128773
rect 232389 128745 232424 128773
rect 232264 128728 232424 128745
rect 247624 128959 247784 128976
rect 247624 128931 247659 128959
rect 247687 128931 247721 128959
rect 247749 128931 247784 128959
rect 247624 128897 247784 128931
rect 247624 128869 247659 128897
rect 247687 128869 247721 128897
rect 247749 128869 247784 128897
rect 247624 128835 247784 128869
rect 247624 128807 247659 128835
rect 247687 128807 247721 128835
rect 247749 128807 247784 128835
rect 247624 128773 247784 128807
rect 247624 128745 247659 128773
rect 247687 128745 247721 128773
rect 247749 128745 247784 128773
rect 247624 128728 247784 128745
rect 254529 128959 254839 137745
rect 254529 128931 254577 128959
rect 254605 128931 254639 128959
rect 254667 128931 254701 128959
rect 254729 128931 254763 128959
rect 254791 128931 254839 128959
rect 254529 128897 254839 128931
rect 254529 128869 254577 128897
rect 254605 128869 254639 128897
rect 254667 128869 254701 128897
rect 254729 128869 254763 128897
rect 254791 128869 254839 128897
rect 254529 128835 254839 128869
rect 254529 128807 254577 128835
rect 254605 128807 254639 128835
rect 254667 128807 254701 128835
rect 254729 128807 254763 128835
rect 254791 128807 254839 128835
rect 254529 128773 254839 128807
rect 254529 128745 254577 128773
rect 254605 128745 254639 128773
rect 254667 128745 254701 128773
rect 254729 128745 254763 128773
rect 254791 128745 254839 128773
rect 31389 122931 31437 122959
rect 31465 122931 31499 122959
rect 31527 122931 31561 122959
rect 31589 122931 31623 122959
rect 31651 122931 31699 122959
rect 31389 122897 31699 122931
rect 31389 122869 31437 122897
rect 31465 122869 31499 122897
rect 31527 122869 31561 122897
rect 31589 122869 31623 122897
rect 31651 122869 31699 122897
rect 31389 122835 31699 122869
rect 31389 122807 31437 122835
rect 31465 122807 31499 122835
rect 31527 122807 31561 122835
rect 31589 122807 31623 122835
rect 31651 122807 31699 122835
rect 31389 122773 31699 122807
rect 31389 122745 31437 122773
rect 31465 122745 31499 122773
rect 31527 122745 31561 122773
rect 31589 122745 31623 122773
rect 31651 122745 31699 122773
rect 31389 113959 31699 122745
rect 40264 122959 40424 122976
rect 40264 122931 40299 122959
rect 40327 122931 40361 122959
rect 40389 122931 40424 122959
rect 40264 122897 40424 122931
rect 40264 122869 40299 122897
rect 40327 122869 40361 122897
rect 40389 122869 40424 122897
rect 40264 122835 40424 122869
rect 40264 122807 40299 122835
rect 40327 122807 40361 122835
rect 40389 122807 40424 122835
rect 40264 122773 40424 122807
rect 40264 122745 40299 122773
rect 40327 122745 40361 122773
rect 40389 122745 40424 122773
rect 40264 122728 40424 122745
rect 55624 122959 55784 122976
rect 55624 122931 55659 122959
rect 55687 122931 55721 122959
rect 55749 122931 55784 122959
rect 55624 122897 55784 122931
rect 55624 122869 55659 122897
rect 55687 122869 55721 122897
rect 55749 122869 55784 122897
rect 55624 122835 55784 122869
rect 55624 122807 55659 122835
rect 55687 122807 55721 122835
rect 55749 122807 55784 122835
rect 55624 122773 55784 122807
rect 55624 122745 55659 122773
rect 55687 122745 55721 122773
rect 55749 122745 55784 122773
rect 55624 122728 55784 122745
rect 70984 122959 71144 122976
rect 70984 122931 71019 122959
rect 71047 122931 71081 122959
rect 71109 122931 71144 122959
rect 70984 122897 71144 122931
rect 70984 122869 71019 122897
rect 71047 122869 71081 122897
rect 71109 122869 71144 122897
rect 70984 122835 71144 122869
rect 70984 122807 71019 122835
rect 71047 122807 71081 122835
rect 71109 122807 71144 122835
rect 70984 122773 71144 122807
rect 70984 122745 71019 122773
rect 71047 122745 71081 122773
rect 71109 122745 71144 122773
rect 70984 122728 71144 122745
rect 86344 122959 86504 122976
rect 86344 122931 86379 122959
rect 86407 122931 86441 122959
rect 86469 122931 86504 122959
rect 86344 122897 86504 122931
rect 86344 122869 86379 122897
rect 86407 122869 86441 122897
rect 86469 122869 86504 122897
rect 86344 122835 86504 122869
rect 86344 122807 86379 122835
rect 86407 122807 86441 122835
rect 86469 122807 86504 122835
rect 86344 122773 86504 122807
rect 86344 122745 86379 122773
rect 86407 122745 86441 122773
rect 86469 122745 86504 122773
rect 86344 122728 86504 122745
rect 101704 122959 101864 122976
rect 101704 122931 101739 122959
rect 101767 122931 101801 122959
rect 101829 122931 101864 122959
rect 101704 122897 101864 122931
rect 101704 122869 101739 122897
rect 101767 122869 101801 122897
rect 101829 122869 101864 122897
rect 101704 122835 101864 122869
rect 101704 122807 101739 122835
rect 101767 122807 101801 122835
rect 101829 122807 101864 122835
rect 101704 122773 101864 122807
rect 101704 122745 101739 122773
rect 101767 122745 101801 122773
rect 101829 122745 101864 122773
rect 101704 122728 101864 122745
rect 117064 122959 117224 122976
rect 117064 122931 117099 122959
rect 117127 122931 117161 122959
rect 117189 122931 117224 122959
rect 117064 122897 117224 122931
rect 117064 122869 117099 122897
rect 117127 122869 117161 122897
rect 117189 122869 117224 122897
rect 117064 122835 117224 122869
rect 117064 122807 117099 122835
rect 117127 122807 117161 122835
rect 117189 122807 117224 122835
rect 117064 122773 117224 122807
rect 117064 122745 117099 122773
rect 117127 122745 117161 122773
rect 117189 122745 117224 122773
rect 117064 122728 117224 122745
rect 132424 122959 132584 122976
rect 132424 122931 132459 122959
rect 132487 122931 132521 122959
rect 132549 122931 132584 122959
rect 132424 122897 132584 122931
rect 132424 122869 132459 122897
rect 132487 122869 132521 122897
rect 132549 122869 132584 122897
rect 132424 122835 132584 122869
rect 132424 122807 132459 122835
rect 132487 122807 132521 122835
rect 132549 122807 132584 122835
rect 132424 122773 132584 122807
rect 132424 122745 132459 122773
rect 132487 122745 132521 122773
rect 132549 122745 132584 122773
rect 132424 122728 132584 122745
rect 147784 122959 147944 122976
rect 147784 122931 147819 122959
rect 147847 122931 147881 122959
rect 147909 122931 147944 122959
rect 147784 122897 147944 122931
rect 147784 122869 147819 122897
rect 147847 122869 147881 122897
rect 147909 122869 147944 122897
rect 147784 122835 147944 122869
rect 147784 122807 147819 122835
rect 147847 122807 147881 122835
rect 147909 122807 147944 122835
rect 147784 122773 147944 122807
rect 147784 122745 147819 122773
rect 147847 122745 147881 122773
rect 147909 122745 147944 122773
rect 147784 122728 147944 122745
rect 163144 122959 163304 122976
rect 163144 122931 163179 122959
rect 163207 122931 163241 122959
rect 163269 122931 163304 122959
rect 163144 122897 163304 122931
rect 163144 122869 163179 122897
rect 163207 122869 163241 122897
rect 163269 122869 163304 122897
rect 163144 122835 163304 122869
rect 163144 122807 163179 122835
rect 163207 122807 163241 122835
rect 163269 122807 163304 122835
rect 163144 122773 163304 122807
rect 163144 122745 163179 122773
rect 163207 122745 163241 122773
rect 163269 122745 163304 122773
rect 163144 122728 163304 122745
rect 178504 122959 178664 122976
rect 178504 122931 178539 122959
rect 178567 122931 178601 122959
rect 178629 122931 178664 122959
rect 178504 122897 178664 122931
rect 178504 122869 178539 122897
rect 178567 122869 178601 122897
rect 178629 122869 178664 122897
rect 178504 122835 178664 122869
rect 178504 122807 178539 122835
rect 178567 122807 178601 122835
rect 178629 122807 178664 122835
rect 178504 122773 178664 122807
rect 178504 122745 178539 122773
rect 178567 122745 178601 122773
rect 178629 122745 178664 122773
rect 178504 122728 178664 122745
rect 193864 122959 194024 122976
rect 193864 122931 193899 122959
rect 193927 122931 193961 122959
rect 193989 122931 194024 122959
rect 193864 122897 194024 122931
rect 193864 122869 193899 122897
rect 193927 122869 193961 122897
rect 193989 122869 194024 122897
rect 193864 122835 194024 122869
rect 193864 122807 193899 122835
rect 193927 122807 193961 122835
rect 193989 122807 194024 122835
rect 193864 122773 194024 122807
rect 193864 122745 193899 122773
rect 193927 122745 193961 122773
rect 193989 122745 194024 122773
rect 193864 122728 194024 122745
rect 209224 122959 209384 122976
rect 209224 122931 209259 122959
rect 209287 122931 209321 122959
rect 209349 122931 209384 122959
rect 209224 122897 209384 122931
rect 209224 122869 209259 122897
rect 209287 122869 209321 122897
rect 209349 122869 209384 122897
rect 209224 122835 209384 122869
rect 209224 122807 209259 122835
rect 209287 122807 209321 122835
rect 209349 122807 209384 122835
rect 209224 122773 209384 122807
rect 209224 122745 209259 122773
rect 209287 122745 209321 122773
rect 209349 122745 209384 122773
rect 209224 122728 209384 122745
rect 224584 122959 224744 122976
rect 224584 122931 224619 122959
rect 224647 122931 224681 122959
rect 224709 122931 224744 122959
rect 224584 122897 224744 122931
rect 224584 122869 224619 122897
rect 224647 122869 224681 122897
rect 224709 122869 224744 122897
rect 224584 122835 224744 122869
rect 224584 122807 224619 122835
rect 224647 122807 224681 122835
rect 224709 122807 224744 122835
rect 224584 122773 224744 122807
rect 224584 122745 224619 122773
rect 224647 122745 224681 122773
rect 224709 122745 224744 122773
rect 224584 122728 224744 122745
rect 239944 122959 240104 122976
rect 239944 122931 239979 122959
rect 240007 122931 240041 122959
rect 240069 122931 240104 122959
rect 239944 122897 240104 122931
rect 239944 122869 239979 122897
rect 240007 122869 240041 122897
rect 240069 122869 240104 122897
rect 239944 122835 240104 122869
rect 239944 122807 239979 122835
rect 240007 122807 240041 122835
rect 240069 122807 240104 122835
rect 239944 122773 240104 122807
rect 239944 122745 239979 122773
rect 240007 122745 240041 122773
rect 240069 122745 240104 122773
rect 239944 122728 240104 122745
rect 32584 119959 32744 119976
rect 32584 119931 32619 119959
rect 32647 119931 32681 119959
rect 32709 119931 32744 119959
rect 32584 119897 32744 119931
rect 32584 119869 32619 119897
rect 32647 119869 32681 119897
rect 32709 119869 32744 119897
rect 32584 119835 32744 119869
rect 32584 119807 32619 119835
rect 32647 119807 32681 119835
rect 32709 119807 32744 119835
rect 32584 119773 32744 119807
rect 32584 119745 32619 119773
rect 32647 119745 32681 119773
rect 32709 119745 32744 119773
rect 32584 119728 32744 119745
rect 47944 119959 48104 119976
rect 47944 119931 47979 119959
rect 48007 119931 48041 119959
rect 48069 119931 48104 119959
rect 47944 119897 48104 119931
rect 47944 119869 47979 119897
rect 48007 119869 48041 119897
rect 48069 119869 48104 119897
rect 47944 119835 48104 119869
rect 47944 119807 47979 119835
rect 48007 119807 48041 119835
rect 48069 119807 48104 119835
rect 47944 119773 48104 119807
rect 47944 119745 47979 119773
rect 48007 119745 48041 119773
rect 48069 119745 48104 119773
rect 47944 119728 48104 119745
rect 63304 119959 63464 119976
rect 63304 119931 63339 119959
rect 63367 119931 63401 119959
rect 63429 119931 63464 119959
rect 63304 119897 63464 119931
rect 63304 119869 63339 119897
rect 63367 119869 63401 119897
rect 63429 119869 63464 119897
rect 63304 119835 63464 119869
rect 63304 119807 63339 119835
rect 63367 119807 63401 119835
rect 63429 119807 63464 119835
rect 63304 119773 63464 119807
rect 63304 119745 63339 119773
rect 63367 119745 63401 119773
rect 63429 119745 63464 119773
rect 63304 119728 63464 119745
rect 78664 119959 78824 119976
rect 78664 119931 78699 119959
rect 78727 119931 78761 119959
rect 78789 119931 78824 119959
rect 78664 119897 78824 119931
rect 78664 119869 78699 119897
rect 78727 119869 78761 119897
rect 78789 119869 78824 119897
rect 78664 119835 78824 119869
rect 78664 119807 78699 119835
rect 78727 119807 78761 119835
rect 78789 119807 78824 119835
rect 78664 119773 78824 119807
rect 78664 119745 78699 119773
rect 78727 119745 78761 119773
rect 78789 119745 78824 119773
rect 78664 119728 78824 119745
rect 94024 119959 94184 119976
rect 94024 119931 94059 119959
rect 94087 119931 94121 119959
rect 94149 119931 94184 119959
rect 94024 119897 94184 119931
rect 94024 119869 94059 119897
rect 94087 119869 94121 119897
rect 94149 119869 94184 119897
rect 94024 119835 94184 119869
rect 94024 119807 94059 119835
rect 94087 119807 94121 119835
rect 94149 119807 94184 119835
rect 94024 119773 94184 119807
rect 94024 119745 94059 119773
rect 94087 119745 94121 119773
rect 94149 119745 94184 119773
rect 94024 119728 94184 119745
rect 109384 119959 109544 119976
rect 109384 119931 109419 119959
rect 109447 119931 109481 119959
rect 109509 119931 109544 119959
rect 109384 119897 109544 119931
rect 109384 119869 109419 119897
rect 109447 119869 109481 119897
rect 109509 119869 109544 119897
rect 109384 119835 109544 119869
rect 109384 119807 109419 119835
rect 109447 119807 109481 119835
rect 109509 119807 109544 119835
rect 109384 119773 109544 119807
rect 109384 119745 109419 119773
rect 109447 119745 109481 119773
rect 109509 119745 109544 119773
rect 109384 119728 109544 119745
rect 124744 119959 124904 119976
rect 124744 119931 124779 119959
rect 124807 119931 124841 119959
rect 124869 119931 124904 119959
rect 124744 119897 124904 119931
rect 124744 119869 124779 119897
rect 124807 119869 124841 119897
rect 124869 119869 124904 119897
rect 124744 119835 124904 119869
rect 124744 119807 124779 119835
rect 124807 119807 124841 119835
rect 124869 119807 124904 119835
rect 124744 119773 124904 119807
rect 124744 119745 124779 119773
rect 124807 119745 124841 119773
rect 124869 119745 124904 119773
rect 124744 119728 124904 119745
rect 140104 119959 140264 119976
rect 140104 119931 140139 119959
rect 140167 119931 140201 119959
rect 140229 119931 140264 119959
rect 140104 119897 140264 119931
rect 140104 119869 140139 119897
rect 140167 119869 140201 119897
rect 140229 119869 140264 119897
rect 140104 119835 140264 119869
rect 140104 119807 140139 119835
rect 140167 119807 140201 119835
rect 140229 119807 140264 119835
rect 140104 119773 140264 119807
rect 140104 119745 140139 119773
rect 140167 119745 140201 119773
rect 140229 119745 140264 119773
rect 140104 119728 140264 119745
rect 155464 119959 155624 119976
rect 155464 119931 155499 119959
rect 155527 119931 155561 119959
rect 155589 119931 155624 119959
rect 155464 119897 155624 119931
rect 155464 119869 155499 119897
rect 155527 119869 155561 119897
rect 155589 119869 155624 119897
rect 155464 119835 155624 119869
rect 155464 119807 155499 119835
rect 155527 119807 155561 119835
rect 155589 119807 155624 119835
rect 155464 119773 155624 119807
rect 155464 119745 155499 119773
rect 155527 119745 155561 119773
rect 155589 119745 155624 119773
rect 155464 119728 155624 119745
rect 170824 119959 170984 119976
rect 170824 119931 170859 119959
rect 170887 119931 170921 119959
rect 170949 119931 170984 119959
rect 170824 119897 170984 119931
rect 170824 119869 170859 119897
rect 170887 119869 170921 119897
rect 170949 119869 170984 119897
rect 170824 119835 170984 119869
rect 170824 119807 170859 119835
rect 170887 119807 170921 119835
rect 170949 119807 170984 119835
rect 170824 119773 170984 119807
rect 170824 119745 170859 119773
rect 170887 119745 170921 119773
rect 170949 119745 170984 119773
rect 170824 119728 170984 119745
rect 186184 119959 186344 119976
rect 186184 119931 186219 119959
rect 186247 119931 186281 119959
rect 186309 119931 186344 119959
rect 186184 119897 186344 119931
rect 186184 119869 186219 119897
rect 186247 119869 186281 119897
rect 186309 119869 186344 119897
rect 186184 119835 186344 119869
rect 186184 119807 186219 119835
rect 186247 119807 186281 119835
rect 186309 119807 186344 119835
rect 186184 119773 186344 119807
rect 186184 119745 186219 119773
rect 186247 119745 186281 119773
rect 186309 119745 186344 119773
rect 186184 119728 186344 119745
rect 201544 119959 201704 119976
rect 201544 119931 201579 119959
rect 201607 119931 201641 119959
rect 201669 119931 201704 119959
rect 201544 119897 201704 119931
rect 201544 119869 201579 119897
rect 201607 119869 201641 119897
rect 201669 119869 201704 119897
rect 201544 119835 201704 119869
rect 201544 119807 201579 119835
rect 201607 119807 201641 119835
rect 201669 119807 201704 119835
rect 201544 119773 201704 119807
rect 201544 119745 201579 119773
rect 201607 119745 201641 119773
rect 201669 119745 201704 119773
rect 201544 119728 201704 119745
rect 216904 119959 217064 119976
rect 216904 119931 216939 119959
rect 216967 119931 217001 119959
rect 217029 119931 217064 119959
rect 216904 119897 217064 119931
rect 216904 119869 216939 119897
rect 216967 119869 217001 119897
rect 217029 119869 217064 119897
rect 216904 119835 217064 119869
rect 216904 119807 216939 119835
rect 216967 119807 217001 119835
rect 217029 119807 217064 119835
rect 216904 119773 217064 119807
rect 216904 119745 216939 119773
rect 216967 119745 217001 119773
rect 217029 119745 217064 119773
rect 216904 119728 217064 119745
rect 232264 119959 232424 119976
rect 232264 119931 232299 119959
rect 232327 119931 232361 119959
rect 232389 119931 232424 119959
rect 232264 119897 232424 119931
rect 232264 119869 232299 119897
rect 232327 119869 232361 119897
rect 232389 119869 232424 119897
rect 232264 119835 232424 119869
rect 232264 119807 232299 119835
rect 232327 119807 232361 119835
rect 232389 119807 232424 119835
rect 232264 119773 232424 119807
rect 232264 119745 232299 119773
rect 232327 119745 232361 119773
rect 232389 119745 232424 119773
rect 232264 119728 232424 119745
rect 247624 119959 247784 119976
rect 247624 119931 247659 119959
rect 247687 119931 247721 119959
rect 247749 119931 247784 119959
rect 247624 119897 247784 119931
rect 247624 119869 247659 119897
rect 247687 119869 247721 119897
rect 247749 119869 247784 119897
rect 247624 119835 247784 119869
rect 247624 119807 247659 119835
rect 247687 119807 247721 119835
rect 247749 119807 247784 119835
rect 247624 119773 247784 119807
rect 247624 119745 247659 119773
rect 247687 119745 247721 119773
rect 247749 119745 247784 119773
rect 247624 119728 247784 119745
rect 254529 119959 254839 128745
rect 254529 119931 254577 119959
rect 254605 119931 254639 119959
rect 254667 119931 254701 119959
rect 254729 119931 254763 119959
rect 254791 119931 254839 119959
rect 254529 119897 254839 119931
rect 254529 119869 254577 119897
rect 254605 119869 254639 119897
rect 254667 119869 254701 119897
rect 254729 119869 254763 119897
rect 254791 119869 254839 119897
rect 254529 119835 254839 119869
rect 254529 119807 254577 119835
rect 254605 119807 254639 119835
rect 254667 119807 254701 119835
rect 254729 119807 254763 119835
rect 254791 119807 254839 119835
rect 254529 119773 254839 119807
rect 254529 119745 254577 119773
rect 254605 119745 254639 119773
rect 254667 119745 254701 119773
rect 254729 119745 254763 119773
rect 254791 119745 254839 119773
rect 31389 113931 31437 113959
rect 31465 113931 31499 113959
rect 31527 113931 31561 113959
rect 31589 113931 31623 113959
rect 31651 113931 31699 113959
rect 31389 113897 31699 113931
rect 31389 113869 31437 113897
rect 31465 113869 31499 113897
rect 31527 113869 31561 113897
rect 31589 113869 31623 113897
rect 31651 113869 31699 113897
rect 31389 113835 31699 113869
rect 31389 113807 31437 113835
rect 31465 113807 31499 113835
rect 31527 113807 31561 113835
rect 31589 113807 31623 113835
rect 31651 113807 31699 113835
rect 31389 113773 31699 113807
rect 31389 113745 31437 113773
rect 31465 113745 31499 113773
rect 31527 113745 31561 113773
rect 31589 113745 31623 113773
rect 31651 113745 31699 113773
rect 31389 104959 31699 113745
rect 40264 113959 40424 113976
rect 40264 113931 40299 113959
rect 40327 113931 40361 113959
rect 40389 113931 40424 113959
rect 40264 113897 40424 113931
rect 40264 113869 40299 113897
rect 40327 113869 40361 113897
rect 40389 113869 40424 113897
rect 40264 113835 40424 113869
rect 40264 113807 40299 113835
rect 40327 113807 40361 113835
rect 40389 113807 40424 113835
rect 40264 113773 40424 113807
rect 40264 113745 40299 113773
rect 40327 113745 40361 113773
rect 40389 113745 40424 113773
rect 40264 113728 40424 113745
rect 55624 113959 55784 113976
rect 55624 113931 55659 113959
rect 55687 113931 55721 113959
rect 55749 113931 55784 113959
rect 55624 113897 55784 113931
rect 55624 113869 55659 113897
rect 55687 113869 55721 113897
rect 55749 113869 55784 113897
rect 55624 113835 55784 113869
rect 55624 113807 55659 113835
rect 55687 113807 55721 113835
rect 55749 113807 55784 113835
rect 55624 113773 55784 113807
rect 55624 113745 55659 113773
rect 55687 113745 55721 113773
rect 55749 113745 55784 113773
rect 55624 113728 55784 113745
rect 70984 113959 71144 113976
rect 70984 113931 71019 113959
rect 71047 113931 71081 113959
rect 71109 113931 71144 113959
rect 70984 113897 71144 113931
rect 70984 113869 71019 113897
rect 71047 113869 71081 113897
rect 71109 113869 71144 113897
rect 70984 113835 71144 113869
rect 70984 113807 71019 113835
rect 71047 113807 71081 113835
rect 71109 113807 71144 113835
rect 70984 113773 71144 113807
rect 70984 113745 71019 113773
rect 71047 113745 71081 113773
rect 71109 113745 71144 113773
rect 70984 113728 71144 113745
rect 86344 113959 86504 113976
rect 86344 113931 86379 113959
rect 86407 113931 86441 113959
rect 86469 113931 86504 113959
rect 86344 113897 86504 113931
rect 86344 113869 86379 113897
rect 86407 113869 86441 113897
rect 86469 113869 86504 113897
rect 86344 113835 86504 113869
rect 86344 113807 86379 113835
rect 86407 113807 86441 113835
rect 86469 113807 86504 113835
rect 86344 113773 86504 113807
rect 86344 113745 86379 113773
rect 86407 113745 86441 113773
rect 86469 113745 86504 113773
rect 86344 113728 86504 113745
rect 101704 113959 101864 113976
rect 101704 113931 101739 113959
rect 101767 113931 101801 113959
rect 101829 113931 101864 113959
rect 101704 113897 101864 113931
rect 101704 113869 101739 113897
rect 101767 113869 101801 113897
rect 101829 113869 101864 113897
rect 101704 113835 101864 113869
rect 101704 113807 101739 113835
rect 101767 113807 101801 113835
rect 101829 113807 101864 113835
rect 101704 113773 101864 113807
rect 101704 113745 101739 113773
rect 101767 113745 101801 113773
rect 101829 113745 101864 113773
rect 101704 113728 101864 113745
rect 117064 113959 117224 113976
rect 117064 113931 117099 113959
rect 117127 113931 117161 113959
rect 117189 113931 117224 113959
rect 117064 113897 117224 113931
rect 117064 113869 117099 113897
rect 117127 113869 117161 113897
rect 117189 113869 117224 113897
rect 117064 113835 117224 113869
rect 117064 113807 117099 113835
rect 117127 113807 117161 113835
rect 117189 113807 117224 113835
rect 117064 113773 117224 113807
rect 117064 113745 117099 113773
rect 117127 113745 117161 113773
rect 117189 113745 117224 113773
rect 117064 113728 117224 113745
rect 132424 113959 132584 113976
rect 132424 113931 132459 113959
rect 132487 113931 132521 113959
rect 132549 113931 132584 113959
rect 132424 113897 132584 113931
rect 132424 113869 132459 113897
rect 132487 113869 132521 113897
rect 132549 113869 132584 113897
rect 132424 113835 132584 113869
rect 132424 113807 132459 113835
rect 132487 113807 132521 113835
rect 132549 113807 132584 113835
rect 132424 113773 132584 113807
rect 132424 113745 132459 113773
rect 132487 113745 132521 113773
rect 132549 113745 132584 113773
rect 132424 113728 132584 113745
rect 147784 113959 147944 113976
rect 147784 113931 147819 113959
rect 147847 113931 147881 113959
rect 147909 113931 147944 113959
rect 147784 113897 147944 113931
rect 147784 113869 147819 113897
rect 147847 113869 147881 113897
rect 147909 113869 147944 113897
rect 147784 113835 147944 113869
rect 147784 113807 147819 113835
rect 147847 113807 147881 113835
rect 147909 113807 147944 113835
rect 147784 113773 147944 113807
rect 147784 113745 147819 113773
rect 147847 113745 147881 113773
rect 147909 113745 147944 113773
rect 147784 113728 147944 113745
rect 163144 113959 163304 113976
rect 163144 113931 163179 113959
rect 163207 113931 163241 113959
rect 163269 113931 163304 113959
rect 163144 113897 163304 113931
rect 163144 113869 163179 113897
rect 163207 113869 163241 113897
rect 163269 113869 163304 113897
rect 163144 113835 163304 113869
rect 163144 113807 163179 113835
rect 163207 113807 163241 113835
rect 163269 113807 163304 113835
rect 163144 113773 163304 113807
rect 163144 113745 163179 113773
rect 163207 113745 163241 113773
rect 163269 113745 163304 113773
rect 163144 113728 163304 113745
rect 178504 113959 178664 113976
rect 178504 113931 178539 113959
rect 178567 113931 178601 113959
rect 178629 113931 178664 113959
rect 178504 113897 178664 113931
rect 178504 113869 178539 113897
rect 178567 113869 178601 113897
rect 178629 113869 178664 113897
rect 178504 113835 178664 113869
rect 178504 113807 178539 113835
rect 178567 113807 178601 113835
rect 178629 113807 178664 113835
rect 178504 113773 178664 113807
rect 178504 113745 178539 113773
rect 178567 113745 178601 113773
rect 178629 113745 178664 113773
rect 178504 113728 178664 113745
rect 193864 113959 194024 113976
rect 193864 113931 193899 113959
rect 193927 113931 193961 113959
rect 193989 113931 194024 113959
rect 193864 113897 194024 113931
rect 193864 113869 193899 113897
rect 193927 113869 193961 113897
rect 193989 113869 194024 113897
rect 193864 113835 194024 113869
rect 193864 113807 193899 113835
rect 193927 113807 193961 113835
rect 193989 113807 194024 113835
rect 193864 113773 194024 113807
rect 193864 113745 193899 113773
rect 193927 113745 193961 113773
rect 193989 113745 194024 113773
rect 193864 113728 194024 113745
rect 209224 113959 209384 113976
rect 209224 113931 209259 113959
rect 209287 113931 209321 113959
rect 209349 113931 209384 113959
rect 209224 113897 209384 113931
rect 209224 113869 209259 113897
rect 209287 113869 209321 113897
rect 209349 113869 209384 113897
rect 209224 113835 209384 113869
rect 209224 113807 209259 113835
rect 209287 113807 209321 113835
rect 209349 113807 209384 113835
rect 209224 113773 209384 113807
rect 209224 113745 209259 113773
rect 209287 113745 209321 113773
rect 209349 113745 209384 113773
rect 209224 113728 209384 113745
rect 224584 113959 224744 113976
rect 224584 113931 224619 113959
rect 224647 113931 224681 113959
rect 224709 113931 224744 113959
rect 224584 113897 224744 113931
rect 224584 113869 224619 113897
rect 224647 113869 224681 113897
rect 224709 113869 224744 113897
rect 224584 113835 224744 113869
rect 224584 113807 224619 113835
rect 224647 113807 224681 113835
rect 224709 113807 224744 113835
rect 224584 113773 224744 113807
rect 224584 113745 224619 113773
rect 224647 113745 224681 113773
rect 224709 113745 224744 113773
rect 224584 113728 224744 113745
rect 239944 113959 240104 113976
rect 239944 113931 239979 113959
rect 240007 113931 240041 113959
rect 240069 113931 240104 113959
rect 239944 113897 240104 113931
rect 239944 113869 239979 113897
rect 240007 113869 240041 113897
rect 240069 113869 240104 113897
rect 239944 113835 240104 113869
rect 239944 113807 239979 113835
rect 240007 113807 240041 113835
rect 240069 113807 240104 113835
rect 239944 113773 240104 113807
rect 239944 113745 239979 113773
rect 240007 113745 240041 113773
rect 240069 113745 240104 113773
rect 239944 113728 240104 113745
rect 32584 110959 32744 110976
rect 32584 110931 32619 110959
rect 32647 110931 32681 110959
rect 32709 110931 32744 110959
rect 32584 110897 32744 110931
rect 32584 110869 32619 110897
rect 32647 110869 32681 110897
rect 32709 110869 32744 110897
rect 32584 110835 32744 110869
rect 32584 110807 32619 110835
rect 32647 110807 32681 110835
rect 32709 110807 32744 110835
rect 32584 110773 32744 110807
rect 32584 110745 32619 110773
rect 32647 110745 32681 110773
rect 32709 110745 32744 110773
rect 32584 110728 32744 110745
rect 47944 110959 48104 110976
rect 47944 110931 47979 110959
rect 48007 110931 48041 110959
rect 48069 110931 48104 110959
rect 47944 110897 48104 110931
rect 47944 110869 47979 110897
rect 48007 110869 48041 110897
rect 48069 110869 48104 110897
rect 47944 110835 48104 110869
rect 47944 110807 47979 110835
rect 48007 110807 48041 110835
rect 48069 110807 48104 110835
rect 47944 110773 48104 110807
rect 47944 110745 47979 110773
rect 48007 110745 48041 110773
rect 48069 110745 48104 110773
rect 47944 110728 48104 110745
rect 63304 110959 63464 110976
rect 63304 110931 63339 110959
rect 63367 110931 63401 110959
rect 63429 110931 63464 110959
rect 63304 110897 63464 110931
rect 63304 110869 63339 110897
rect 63367 110869 63401 110897
rect 63429 110869 63464 110897
rect 63304 110835 63464 110869
rect 63304 110807 63339 110835
rect 63367 110807 63401 110835
rect 63429 110807 63464 110835
rect 63304 110773 63464 110807
rect 63304 110745 63339 110773
rect 63367 110745 63401 110773
rect 63429 110745 63464 110773
rect 63304 110728 63464 110745
rect 78664 110959 78824 110976
rect 78664 110931 78699 110959
rect 78727 110931 78761 110959
rect 78789 110931 78824 110959
rect 78664 110897 78824 110931
rect 78664 110869 78699 110897
rect 78727 110869 78761 110897
rect 78789 110869 78824 110897
rect 78664 110835 78824 110869
rect 78664 110807 78699 110835
rect 78727 110807 78761 110835
rect 78789 110807 78824 110835
rect 78664 110773 78824 110807
rect 78664 110745 78699 110773
rect 78727 110745 78761 110773
rect 78789 110745 78824 110773
rect 78664 110728 78824 110745
rect 94024 110959 94184 110976
rect 94024 110931 94059 110959
rect 94087 110931 94121 110959
rect 94149 110931 94184 110959
rect 94024 110897 94184 110931
rect 94024 110869 94059 110897
rect 94087 110869 94121 110897
rect 94149 110869 94184 110897
rect 94024 110835 94184 110869
rect 94024 110807 94059 110835
rect 94087 110807 94121 110835
rect 94149 110807 94184 110835
rect 94024 110773 94184 110807
rect 94024 110745 94059 110773
rect 94087 110745 94121 110773
rect 94149 110745 94184 110773
rect 94024 110728 94184 110745
rect 109384 110959 109544 110976
rect 109384 110931 109419 110959
rect 109447 110931 109481 110959
rect 109509 110931 109544 110959
rect 109384 110897 109544 110931
rect 109384 110869 109419 110897
rect 109447 110869 109481 110897
rect 109509 110869 109544 110897
rect 109384 110835 109544 110869
rect 109384 110807 109419 110835
rect 109447 110807 109481 110835
rect 109509 110807 109544 110835
rect 109384 110773 109544 110807
rect 109384 110745 109419 110773
rect 109447 110745 109481 110773
rect 109509 110745 109544 110773
rect 109384 110728 109544 110745
rect 124744 110959 124904 110976
rect 124744 110931 124779 110959
rect 124807 110931 124841 110959
rect 124869 110931 124904 110959
rect 124744 110897 124904 110931
rect 124744 110869 124779 110897
rect 124807 110869 124841 110897
rect 124869 110869 124904 110897
rect 124744 110835 124904 110869
rect 124744 110807 124779 110835
rect 124807 110807 124841 110835
rect 124869 110807 124904 110835
rect 124744 110773 124904 110807
rect 124744 110745 124779 110773
rect 124807 110745 124841 110773
rect 124869 110745 124904 110773
rect 124744 110728 124904 110745
rect 140104 110959 140264 110976
rect 140104 110931 140139 110959
rect 140167 110931 140201 110959
rect 140229 110931 140264 110959
rect 140104 110897 140264 110931
rect 140104 110869 140139 110897
rect 140167 110869 140201 110897
rect 140229 110869 140264 110897
rect 140104 110835 140264 110869
rect 140104 110807 140139 110835
rect 140167 110807 140201 110835
rect 140229 110807 140264 110835
rect 140104 110773 140264 110807
rect 140104 110745 140139 110773
rect 140167 110745 140201 110773
rect 140229 110745 140264 110773
rect 140104 110728 140264 110745
rect 155464 110959 155624 110976
rect 155464 110931 155499 110959
rect 155527 110931 155561 110959
rect 155589 110931 155624 110959
rect 155464 110897 155624 110931
rect 155464 110869 155499 110897
rect 155527 110869 155561 110897
rect 155589 110869 155624 110897
rect 155464 110835 155624 110869
rect 155464 110807 155499 110835
rect 155527 110807 155561 110835
rect 155589 110807 155624 110835
rect 155464 110773 155624 110807
rect 155464 110745 155499 110773
rect 155527 110745 155561 110773
rect 155589 110745 155624 110773
rect 155464 110728 155624 110745
rect 170824 110959 170984 110976
rect 170824 110931 170859 110959
rect 170887 110931 170921 110959
rect 170949 110931 170984 110959
rect 170824 110897 170984 110931
rect 170824 110869 170859 110897
rect 170887 110869 170921 110897
rect 170949 110869 170984 110897
rect 170824 110835 170984 110869
rect 170824 110807 170859 110835
rect 170887 110807 170921 110835
rect 170949 110807 170984 110835
rect 170824 110773 170984 110807
rect 170824 110745 170859 110773
rect 170887 110745 170921 110773
rect 170949 110745 170984 110773
rect 170824 110728 170984 110745
rect 186184 110959 186344 110976
rect 186184 110931 186219 110959
rect 186247 110931 186281 110959
rect 186309 110931 186344 110959
rect 186184 110897 186344 110931
rect 186184 110869 186219 110897
rect 186247 110869 186281 110897
rect 186309 110869 186344 110897
rect 186184 110835 186344 110869
rect 186184 110807 186219 110835
rect 186247 110807 186281 110835
rect 186309 110807 186344 110835
rect 186184 110773 186344 110807
rect 186184 110745 186219 110773
rect 186247 110745 186281 110773
rect 186309 110745 186344 110773
rect 186184 110728 186344 110745
rect 201544 110959 201704 110976
rect 201544 110931 201579 110959
rect 201607 110931 201641 110959
rect 201669 110931 201704 110959
rect 201544 110897 201704 110931
rect 201544 110869 201579 110897
rect 201607 110869 201641 110897
rect 201669 110869 201704 110897
rect 201544 110835 201704 110869
rect 201544 110807 201579 110835
rect 201607 110807 201641 110835
rect 201669 110807 201704 110835
rect 201544 110773 201704 110807
rect 201544 110745 201579 110773
rect 201607 110745 201641 110773
rect 201669 110745 201704 110773
rect 201544 110728 201704 110745
rect 216904 110959 217064 110976
rect 216904 110931 216939 110959
rect 216967 110931 217001 110959
rect 217029 110931 217064 110959
rect 216904 110897 217064 110931
rect 216904 110869 216939 110897
rect 216967 110869 217001 110897
rect 217029 110869 217064 110897
rect 216904 110835 217064 110869
rect 216904 110807 216939 110835
rect 216967 110807 217001 110835
rect 217029 110807 217064 110835
rect 216904 110773 217064 110807
rect 216904 110745 216939 110773
rect 216967 110745 217001 110773
rect 217029 110745 217064 110773
rect 216904 110728 217064 110745
rect 232264 110959 232424 110976
rect 232264 110931 232299 110959
rect 232327 110931 232361 110959
rect 232389 110931 232424 110959
rect 232264 110897 232424 110931
rect 232264 110869 232299 110897
rect 232327 110869 232361 110897
rect 232389 110869 232424 110897
rect 232264 110835 232424 110869
rect 232264 110807 232299 110835
rect 232327 110807 232361 110835
rect 232389 110807 232424 110835
rect 232264 110773 232424 110807
rect 232264 110745 232299 110773
rect 232327 110745 232361 110773
rect 232389 110745 232424 110773
rect 232264 110728 232424 110745
rect 247624 110959 247784 110976
rect 247624 110931 247659 110959
rect 247687 110931 247721 110959
rect 247749 110931 247784 110959
rect 247624 110897 247784 110931
rect 247624 110869 247659 110897
rect 247687 110869 247721 110897
rect 247749 110869 247784 110897
rect 247624 110835 247784 110869
rect 247624 110807 247659 110835
rect 247687 110807 247721 110835
rect 247749 110807 247784 110835
rect 247624 110773 247784 110807
rect 247624 110745 247659 110773
rect 247687 110745 247721 110773
rect 247749 110745 247784 110773
rect 247624 110728 247784 110745
rect 254529 110959 254839 119745
rect 254529 110931 254577 110959
rect 254605 110931 254639 110959
rect 254667 110931 254701 110959
rect 254729 110931 254763 110959
rect 254791 110931 254839 110959
rect 254529 110897 254839 110931
rect 254529 110869 254577 110897
rect 254605 110869 254639 110897
rect 254667 110869 254701 110897
rect 254729 110869 254763 110897
rect 254791 110869 254839 110897
rect 254529 110835 254839 110869
rect 254529 110807 254577 110835
rect 254605 110807 254639 110835
rect 254667 110807 254701 110835
rect 254729 110807 254763 110835
rect 254791 110807 254839 110835
rect 254529 110773 254839 110807
rect 254529 110745 254577 110773
rect 254605 110745 254639 110773
rect 254667 110745 254701 110773
rect 254729 110745 254763 110773
rect 254791 110745 254839 110773
rect 31389 104931 31437 104959
rect 31465 104931 31499 104959
rect 31527 104931 31561 104959
rect 31589 104931 31623 104959
rect 31651 104931 31699 104959
rect 31389 104897 31699 104931
rect 31389 104869 31437 104897
rect 31465 104869 31499 104897
rect 31527 104869 31561 104897
rect 31589 104869 31623 104897
rect 31651 104869 31699 104897
rect 31389 104835 31699 104869
rect 31389 104807 31437 104835
rect 31465 104807 31499 104835
rect 31527 104807 31561 104835
rect 31589 104807 31623 104835
rect 31651 104807 31699 104835
rect 31389 104773 31699 104807
rect 31389 104745 31437 104773
rect 31465 104745 31499 104773
rect 31527 104745 31561 104773
rect 31589 104745 31623 104773
rect 31651 104745 31699 104773
rect 31389 95959 31699 104745
rect 40264 104959 40424 104976
rect 40264 104931 40299 104959
rect 40327 104931 40361 104959
rect 40389 104931 40424 104959
rect 40264 104897 40424 104931
rect 40264 104869 40299 104897
rect 40327 104869 40361 104897
rect 40389 104869 40424 104897
rect 40264 104835 40424 104869
rect 40264 104807 40299 104835
rect 40327 104807 40361 104835
rect 40389 104807 40424 104835
rect 40264 104773 40424 104807
rect 40264 104745 40299 104773
rect 40327 104745 40361 104773
rect 40389 104745 40424 104773
rect 40264 104728 40424 104745
rect 55624 104959 55784 104976
rect 55624 104931 55659 104959
rect 55687 104931 55721 104959
rect 55749 104931 55784 104959
rect 55624 104897 55784 104931
rect 55624 104869 55659 104897
rect 55687 104869 55721 104897
rect 55749 104869 55784 104897
rect 55624 104835 55784 104869
rect 55624 104807 55659 104835
rect 55687 104807 55721 104835
rect 55749 104807 55784 104835
rect 55624 104773 55784 104807
rect 55624 104745 55659 104773
rect 55687 104745 55721 104773
rect 55749 104745 55784 104773
rect 55624 104728 55784 104745
rect 70984 104959 71144 104976
rect 70984 104931 71019 104959
rect 71047 104931 71081 104959
rect 71109 104931 71144 104959
rect 70984 104897 71144 104931
rect 70984 104869 71019 104897
rect 71047 104869 71081 104897
rect 71109 104869 71144 104897
rect 70984 104835 71144 104869
rect 70984 104807 71019 104835
rect 71047 104807 71081 104835
rect 71109 104807 71144 104835
rect 70984 104773 71144 104807
rect 70984 104745 71019 104773
rect 71047 104745 71081 104773
rect 71109 104745 71144 104773
rect 70984 104728 71144 104745
rect 86344 104959 86504 104976
rect 86344 104931 86379 104959
rect 86407 104931 86441 104959
rect 86469 104931 86504 104959
rect 86344 104897 86504 104931
rect 86344 104869 86379 104897
rect 86407 104869 86441 104897
rect 86469 104869 86504 104897
rect 86344 104835 86504 104869
rect 86344 104807 86379 104835
rect 86407 104807 86441 104835
rect 86469 104807 86504 104835
rect 86344 104773 86504 104807
rect 86344 104745 86379 104773
rect 86407 104745 86441 104773
rect 86469 104745 86504 104773
rect 86344 104728 86504 104745
rect 101704 104959 101864 104976
rect 101704 104931 101739 104959
rect 101767 104931 101801 104959
rect 101829 104931 101864 104959
rect 101704 104897 101864 104931
rect 101704 104869 101739 104897
rect 101767 104869 101801 104897
rect 101829 104869 101864 104897
rect 101704 104835 101864 104869
rect 101704 104807 101739 104835
rect 101767 104807 101801 104835
rect 101829 104807 101864 104835
rect 101704 104773 101864 104807
rect 101704 104745 101739 104773
rect 101767 104745 101801 104773
rect 101829 104745 101864 104773
rect 101704 104728 101864 104745
rect 117064 104959 117224 104976
rect 117064 104931 117099 104959
rect 117127 104931 117161 104959
rect 117189 104931 117224 104959
rect 117064 104897 117224 104931
rect 117064 104869 117099 104897
rect 117127 104869 117161 104897
rect 117189 104869 117224 104897
rect 117064 104835 117224 104869
rect 117064 104807 117099 104835
rect 117127 104807 117161 104835
rect 117189 104807 117224 104835
rect 117064 104773 117224 104807
rect 117064 104745 117099 104773
rect 117127 104745 117161 104773
rect 117189 104745 117224 104773
rect 117064 104728 117224 104745
rect 132424 104959 132584 104976
rect 132424 104931 132459 104959
rect 132487 104931 132521 104959
rect 132549 104931 132584 104959
rect 132424 104897 132584 104931
rect 132424 104869 132459 104897
rect 132487 104869 132521 104897
rect 132549 104869 132584 104897
rect 132424 104835 132584 104869
rect 132424 104807 132459 104835
rect 132487 104807 132521 104835
rect 132549 104807 132584 104835
rect 132424 104773 132584 104807
rect 132424 104745 132459 104773
rect 132487 104745 132521 104773
rect 132549 104745 132584 104773
rect 132424 104728 132584 104745
rect 147784 104959 147944 104976
rect 147784 104931 147819 104959
rect 147847 104931 147881 104959
rect 147909 104931 147944 104959
rect 147784 104897 147944 104931
rect 147784 104869 147819 104897
rect 147847 104869 147881 104897
rect 147909 104869 147944 104897
rect 147784 104835 147944 104869
rect 147784 104807 147819 104835
rect 147847 104807 147881 104835
rect 147909 104807 147944 104835
rect 147784 104773 147944 104807
rect 147784 104745 147819 104773
rect 147847 104745 147881 104773
rect 147909 104745 147944 104773
rect 147784 104728 147944 104745
rect 163144 104959 163304 104976
rect 163144 104931 163179 104959
rect 163207 104931 163241 104959
rect 163269 104931 163304 104959
rect 163144 104897 163304 104931
rect 163144 104869 163179 104897
rect 163207 104869 163241 104897
rect 163269 104869 163304 104897
rect 163144 104835 163304 104869
rect 163144 104807 163179 104835
rect 163207 104807 163241 104835
rect 163269 104807 163304 104835
rect 163144 104773 163304 104807
rect 163144 104745 163179 104773
rect 163207 104745 163241 104773
rect 163269 104745 163304 104773
rect 163144 104728 163304 104745
rect 178504 104959 178664 104976
rect 178504 104931 178539 104959
rect 178567 104931 178601 104959
rect 178629 104931 178664 104959
rect 178504 104897 178664 104931
rect 178504 104869 178539 104897
rect 178567 104869 178601 104897
rect 178629 104869 178664 104897
rect 178504 104835 178664 104869
rect 178504 104807 178539 104835
rect 178567 104807 178601 104835
rect 178629 104807 178664 104835
rect 178504 104773 178664 104807
rect 178504 104745 178539 104773
rect 178567 104745 178601 104773
rect 178629 104745 178664 104773
rect 178504 104728 178664 104745
rect 193864 104959 194024 104976
rect 193864 104931 193899 104959
rect 193927 104931 193961 104959
rect 193989 104931 194024 104959
rect 193864 104897 194024 104931
rect 193864 104869 193899 104897
rect 193927 104869 193961 104897
rect 193989 104869 194024 104897
rect 193864 104835 194024 104869
rect 193864 104807 193899 104835
rect 193927 104807 193961 104835
rect 193989 104807 194024 104835
rect 193864 104773 194024 104807
rect 193864 104745 193899 104773
rect 193927 104745 193961 104773
rect 193989 104745 194024 104773
rect 193864 104728 194024 104745
rect 209224 104959 209384 104976
rect 209224 104931 209259 104959
rect 209287 104931 209321 104959
rect 209349 104931 209384 104959
rect 209224 104897 209384 104931
rect 209224 104869 209259 104897
rect 209287 104869 209321 104897
rect 209349 104869 209384 104897
rect 209224 104835 209384 104869
rect 209224 104807 209259 104835
rect 209287 104807 209321 104835
rect 209349 104807 209384 104835
rect 209224 104773 209384 104807
rect 209224 104745 209259 104773
rect 209287 104745 209321 104773
rect 209349 104745 209384 104773
rect 209224 104728 209384 104745
rect 224584 104959 224744 104976
rect 224584 104931 224619 104959
rect 224647 104931 224681 104959
rect 224709 104931 224744 104959
rect 224584 104897 224744 104931
rect 224584 104869 224619 104897
rect 224647 104869 224681 104897
rect 224709 104869 224744 104897
rect 224584 104835 224744 104869
rect 224584 104807 224619 104835
rect 224647 104807 224681 104835
rect 224709 104807 224744 104835
rect 224584 104773 224744 104807
rect 224584 104745 224619 104773
rect 224647 104745 224681 104773
rect 224709 104745 224744 104773
rect 224584 104728 224744 104745
rect 239944 104959 240104 104976
rect 239944 104931 239979 104959
rect 240007 104931 240041 104959
rect 240069 104931 240104 104959
rect 239944 104897 240104 104931
rect 239944 104869 239979 104897
rect 240007 104869 240041 104897
rect 240069 104869 240104 104897
rect 239944 104835 240104 104869
rect 239944 104807 239979 104835
rect 240007 104807 240041 104835
rect 240069 104807 240104 104835
rect 239944 104773 240104 104807
rect 239944 104745 239979 104773
rect 240007 104745 240041 104773
rect 240069 104745 240104 104773
rect 239944 104728 240104 104745
rect 32584 101959 32744 101976
rect 32584 101931 32619 101959
rect 32647 101931 32681 101959
rect 32709 101931 32744 101959
rect 32584 101897 32744 101931
rect 32584 101869 32619 101897
rect 32647 101869 32681 101897
rect 32709 101869 32744 101897
rect 32584 101835 32744 101869
rect 32584 101807 32619 101835
rect 32647 101807 32681 101835
rect 32709 101807 32744 101835
rect 32584 101773 32744 101807
rect 32584 101745 32619 101773
rect 32647 101745 32681 101773
rect 32709 101745 32744 101773
rect 32584 101728 32744 101745
rect 47944 101959 48104 101976
rect 47944 101931 47979 101959
rect 48007 101931 48041 101959
rect 48069 101931 48104 101959
rect 47944 101897 48104 101931
rect 47944 101869 47979 101897
rect 48007 101869 48041 101897
rect 48069 101869 48104 101897
rect 47944 101835 48104 101869
rect 47944 101807 47979 101835
rect 48007 101807 48041 101835
rect 48069 101807 48104 101835
rect 47944 101773 48104 101807
rect 47944 101745 47979 101773
rect 48007 101745 48041 101773
rect 48069 101745 48104 101773
rect 47944 101728 48104 101745
rect 63304 101959 63464 101976
rect 63304 101931 63339 101959
rect 63367 101931 63401 101959
rect 63429 101931 63464 101959
rect 63304 101897 63464 101931
rect 63304 101869 63339 101897
rect 63367 101869 63401 101897
rect 63429 101869 63464 101897
rect 63304 101835 63464 101869
rect 63304 101807 63339 101835
rect 63367 101807 63401 101835
rect 63429 101807 63464 101835
rect 63304 101773 63464 101807
rect 63304 101745 63339 101773
rect 63367 101745 63401 101773
rect 63429 101745 63464 101773
rect 63304 101728 63464 101745
rect 78664 101959 78824 101976
rect 78664 101931 78699 101959
rect 78727 101931 78761 101959
rect 78789 101931 78824 101959
rect 78664 101897 78824 101931
rect 78664 101869 78699 101897
rect 78727 101869 78761 101897
rect 78789 101869 78824 101897
rect 78664 101835 78824 101869
rect 78664 101807 78699 101835
rect 78727 101807 78761 101835
rect 78789 101807 78824 101835
rect 78664 101773 78824 101807
rect 78664 101745 78699 101773
rect 78727 101745 78761 101773
rect 78789 101745 78824 101773
rect 78664 101728 78824 101745
rect 94024 101959 94184 101976
rect 94024 101931 94059 101959
rect 94087 101931 94121 101959
rect 94149 101931 94184 101959
rect 94024 101897 94184 101931
rect 94024 101869 94059 101897
rect 94087 101869 94121 101897
rect 94149 101869 94184 101897
rect 94024 101835 94184 101869
rect 94024 101807 94059 101835
rect 94087 101807 94121 101835
rect 94149 101807 94184 101835
rect 94024 101773 94184 101807
rect 94024 101745 94059 101773
rect 94087 101745 94121 101773
rect 94149 101745 94184 101773
rect 94024 101728 94184 101745
rect 109384 101959 109544 101976
rect 109384 101931 109419 101959
rect 109447 101931 109481 101959
rect 109509 101931 109544 101959
rect 109384 101897 109544 101931
rect 109384 101869 109419 101897
rect 109447 101869 109481 101897
rect 109509 101869 109544 101897
rect 109384 101835 109544 101869
rect 109384 101807 109419 101835
rect 109447 101807 109481 101835
rect 109509 101807 109544 101835
rect 109384 101773 109544 101807
rect 109384 101745 109419 101773
rect 109447 101745 109481 101773
rect 109509 101745 109544 101773
rect 109384 101728 109544 101745
rect 124744 101959 124904 101976
rect 124744 101931 124779 101959
rect 124807 101931 124841 101959
rect 124869 101931 124904 101959
rect 124744 101897 124904 101931
rect 124744 101869 124779 101897
rect 124807 101869 124841 101897
rect 124869 101869 124904 101897
rect 124744 101835 124904 101869
rect 124744 101807 124779 101835
rect 124807 101807 124841 101835
rect 124869 101807 124904 101835
rect 124744 101773 124904 101807
rect 124744 101745 124779 101773
rect 124807 101745 124841 101773
rect 124869 101745 124904 101773
rect 124744 101728 124904 101745
rect 140104 101959 140264 101976
rect 140104 101931 140139 101959
rect 140167 101931 140201 101959
rect 140229 101931 140264 101959
rect 140104 101897 140264 101931
rect 140104 101869 140139 101897
rect 140167 101869 140201 101897
rect 140229 101869 140264 101897
rect 140104 101835 140264 101869
rect 140104 101807 140139 101835
rect 140167 101807 140201 101835
rect 140229 101807 140264 101835
rect 140104 101773 140264 101807
rect 140104 101745 140139 101773
rect 140167 101745 140201 101773
rect 140229 101745 140264 101773
rect 140104 101728 140264 101745
rect 155464 101959 155624 101976
rect 155464 101931 155499 101959
rect 155527 101931 155561 101959
rect 155589 101931 155624 101959
rect 155464 101897 155624 101931
rect 155464 101869 155499 101897
rect 155527 101869 155561 101897
rect 155589 101869 155624 101897
rect 155464 101835 155624 101869
rect 155464 101807 155499 101835
rect 155527 101807 155561 101835
rect 155589 101807 155624 101835
rect 155464 101773 155624 101807
rect 155464 101745 155499 101773
rect 155527 101745 155561 101773
rect 155589 101745 155624 101773
rect 155464 101728 155624 101745
rect 170824 101959 170984 101976
rect 170824 101931 170859 101959
rect 170887 101931 170921 101959
rect 170949 101931 170984 101959
rect 170824 101897 170984 101931
rect 170824 101869 170859 101897
rect 170887 101869 170921 101897
rect 170949 101869 170984 101897
rect 170824 101835 170984 101869
rect 170824 101807 170859 101835
rect 170887 101807 170921 101835
rect 170949 101807 170984 101835
rect 170824 101773 170984 101807
rect 170824 101745 170859 101773
rect 170887 101745 170921 101773
rect 170949 101745 170984 101773
rect 170824 101728 170984 101745
rect 186184 101959 186344 101976
rect 186184 101931 186219 101959
rect 186247 101931 186281 101959
rect 186309 101931 186344 101959
rect 186184 101897 186344 101931
rect 186184 101869 186219 101897
rect 186247 101869 186281 101897
rect 186309 101869 186344 101897
rect 186184 101835 186344 101869
rect 186184 101807 186219 101835
rect 186247 101807 186281 101835
rect 186309 101807 186344 101835
rect 186184 101773 186344 101807
rect 186184 101745 186219 101773
rect 186247 101745 186281 101773
rect 186309 101745 186344 101773
rect 186184 101728 186344 101745
rect 201544 101959 201704 101976
rect 201544 101931 201579 101959
rect 201607 101931 201641 101959
rect 201669 101931 201704 101959
rect 201544 101897 201704 101931
rect 201544 101869 201579 101897
rect 201607 101869 201641 101897
rect 201669 101869 201704 101897
rect 201544 101835 201704 101869
rect 201544 101807 201579 101835
rect 201607 101807 201641 101835
rect 201669 101807 201704 101835
rect 201544 101773 201704 101807
rect 201544 101745 201579 101773
rect 201607 101745 201641 101773
rect 201669 101745 201704 101773
rect 201544 101728 201704 101745
rect 216904 101959 217064 101976
rect 216904 101931 216939 101959
rect 216967 101931 217001 101959
rect 217029 101931 217064 101959
rect 216904 101897 217064 101931
rect 216904 101869 216939 101897
rect 216967 101869 217001 101897
rect 217029 101869 217064 101897
rect 216904 101835 217064 101869
rect 216904 101807 216939 101835
rect 216967 101807 217001 101835
rect 217029 101807 217064 101835
rect 216904 101773 217064 101807
rect 216904 101745 216939 101773
rect 216967 101745 217001 101773
rect 217029 101745 217064 101773
rect 216904 101728 217064 101745
rect 232264 101959 232424 101976
rect 232264 101931 232299 101959
rect 232327 101931 232361 101959
rect 232389 101931 232424 101959
rect 232264 101897 232424 101931
rect 232264 101869 232299 101897
rect 232327 101869 232361 101897
rect 232389 101869 232424 101897
rect 232264 101835 232424 101869
rect 232264 101807 232299 101835
rect 232327 101807 232361 101835
rect 232389 101807 232424 101835
rect 232264 101773 232424 101807
rect 232264 101745 232299 101773
rect 232327 101745 232361 101773
rect 232389 101745 232424 101773
rect 232264 101728 232424 101745
rect 247624 101959 247784 101976
rect 247624 101931 247659 101959
rect 247687 101931 247721 101959
rect 247749 101931 247784 101959
rect 247624 101897 247784 101931
rect 247624 101869 247659 101897
rect 247687 101869 247721 101897
rect 247749 101869 247784 101897
rect 247624 101835 247784 101869
rect 247624 101807 247659 101835
rect 247687 101807 247721 101835
rect 247749 101807 247784 101835
rect 247624 101773 247784 101807
rect 247624 101745 247659 101773
rect 247687 101745 247721 101773
rect 247749 101745 247784 101773
rect 247624 101728 247784 101745
rect 254529 101959 254839 110745
rect 254529 101931 254577 101959
rect 254605 101931 254639 101959
rect 254667 101931 254701 101959
rect 254729 101931 254763 101959
rect 254791 101931 254839 101959
rect 254529 101897 254839 101931
rect 254529 101869 254577 101897
rect 254605 101869 254639 101897
rect 254667 101869 254701 101897
rect 254729 101869 254763 101897
rect 254791 101869 254839 101897
rect 254529 101835 254839 101869
rect 254529 101807 254577 101835
rect 254605 101807 254639 101835
rect 254667 101807 254701 101835
rect 254729 101807 254763 101835
rect 254791 101807 254839 101835
rect 254529 101773 254839 101807
rect 254529 101745 254577 101773
rect 254605 101745 254639 101773
rect 254667 101745 254701 101773
rect 254729 101745 254763 101773
rect 254791 101745 254839 101773
rect 31389 95931 31437 95959
rect 31465 95931 31499 95959
rect 31527 95931 31561 95959
rect 31589 95931 31623 95959
rect 31651 95931 31699 95959
rect 31389 95897 31699 95931
rect 31389 95869 31437 95897
rect 31465 95869 31499 95897
rect 31527 95869 31561 95897
rect 31589 95869 31623 95897
rect 31651 95869 31699 95897
rect 31389 95835 31699 95869
rect 31389 95807 31437 95835
rect 31465 95807 31499 95835
rect 31527 95807 31561 95835
rect 31589 95807 31623 95835
rect 31651 95807 31699 95835
rect 31389 95773 31699 95807
rect 31389 95745 31437 95773
rect 31465 95745 31499 95773
rect 31527 95745 31561 95773
rect 31589 95745 31623 95773
rect 31651 95745 31699 95773
rect 31389 86959 31699 95745
rect 40264 95959 40424 95976
rect 40264 95931 40299 95959
rect 40327 95931 40361 95959
rect 40389 95931 40424 95959
rect 40264 95897 40424 95931
rect 40264 95869 40299 95897
rect 40327 95869 40361 95897
rect 40389 95869 40424 95897
rect 40264 95835 40424 95869
rect 40264 95807 40299 95835
rect 40327 95807 40361 95835
rect 40389 95807 40424 95835
rect 40264 95773 40424 95807
rect 40264 95745 40299 95773
rect 40327 95745 40361 95773
rect 40389 95745 40424 95773
rect 40264 95728 40424 95745
rect 55624 95959 55784 95976
rect 55624 95931 55659 95959
rect 55687 95931 55721 95959
rect 55749 95931 55784 95959
rect 55624 95897 55784 95931
rect 55624 95869 55659 95897
rect 55687 95869 55721 95897
rect 55749 95869 55784 95897
rect 55624 95835 55784 95869
rect 55624 95807 55659 95835
rect 55687 95807 55721 95835
rect 55749 95807 55784 95835
rect 55624 95773 55784 95807
rect 55624 95745 55659 95773
rect 55687 95745 55721 95773
rect 55749 95745 55784 95773
rect 55624 95728 55784 95745
rect 70984 95959 71144 95976
rect 70984 95931 71019 95959
rect 71047 95931 71081 95959
rect 71109 95931 71144 95959
rect 70984 95897 71144 95931
rect 70984 95869 71019 95897
rect 71047 95869 71081 95897
rect 71109 95869 71144 95897
rect 70984 95835 71144 95869
rect 70984 95807 71019 95835
rect 71047 95807 71081 95835
rect 71109 95807 71144 95835
rect 70984 95773 71144 95807
rect 70984 95745 71019 95773
rect 71047 95745 71081 95773
rect 71109 95745 71144 95773
rect 70984 95728 71144 95745
rect 86344 95959 86504 95976
rect 86344 95931 86379 95959
rect 86407 95931 86441 95959
rect 86469 95931 86504 95959
rect 86344 95897 86504 95931
rect 86344 95869 86379 95897
rect 86407 95869 86441 95897
rect 86469 95869 86504 95897
rect 86344 95835 86504 95869
rect 86344 95807 86379 95835
rect 86407 95807 86441 95835
rect 86469 95807 86504 95835
rect 86344 95773 86504 95807
rect 86344 95745 86379 95773
rect 86407 95745 86441 95773
rect 86469 95745 86504 95773
rect 86344 95728 86504 95745
rect 101704 95959 101864 95976
rect 101704 95931 101739 95959
rect 101767 95931 101801 95959
rect 101829 95931 101864 95959
rect 101704 95897 101864 95931
rect 101704 95869 101739 95897
rect 101767 95869 101801 95897
rect 101829 95869 101864 95897
rect 101704 95835 101864 95869
rect 101704 95807 101739 95835
rect 101767 95807 101801 95835
rect 101829 95807 101864 95835
rect 101704 95773 101864 95807
rect 101704 95745 101739 95773
rect 101767 95745 101801 95773
rect 101829 95745 101864 95773
rect 101704 95728 101864 95745
rect 117064 95959 117224 95976
rect 117064 95931 117099 95959
rect 117127 95931 117161 95959
rect 117189 95931 117224 95959
rect 117064 95897 117224 95931
rect 117064 95869 117099 95897
rect 117127 95869 117161 95897
rect 117189 95869 117224 95897
rect 117064 95835 117224 95869
rect 117064 95807 117099 95835
rect 117127 95807 117161 95835
rect 117189 95807 117224 95835
rect 117064 95773 117224 95807
rect 117064 95745 117099 95773
rect 117127 95745 117161 95773
rect 117189 95745 117224 95773
rect 117064 95728 117224 95745
rect 132424 95959 132584 95976
rect 132424 95931 132459 95959
rect 132487 95931 132521 95959
rect 132549 95931 132584 95959
rect 132424 95897 132584 95931
rect 132424 95869 132459 95897
rect 132487 95869 132521 95897
rect 132549 95869 132584 95897
rect 132424 95835 132584 95869
rect 132424 95807 132459 95835
rect 132487 95807 132521 95835
rect 132549 95807 132584 95835
rect 132424 95773 132584 95807
rect 132424 95745 132459 95773
rect 132487 95745 132521 95773
rect 132549 95745 132584 95773
rect 132424 95728 132584 95745
rect 147784 95959 147944 95976
rect 147784 95931 147819 95959
rect 147847 95931 147881 95959
rect 147909 95931 147944 95959
rect 147784 95897 147944 95931
rect 147784 95869 147819 95897
rect 147847 95869 147881 95897
rect 147909 95869 147944 95897
rect 147784 95835 147944 95869
rect 147784 95807 147819 95835
rect 147847 95807 147881 95835
rect 147909 95807 147944 95835
rect 147784 95773 147944 95807
rect 147784 95745 147819 95773
rect 147847 95745 147881 95773
rect 147909 95745 147944 95773
rect 147784 95728 147944 95745
rect 163144 95959 163304 95976
rect 163144 95931 163179 95959
rect 163207 95931 163241 95959
rect 163269 95931 163304 95959
rect 163144 95897 163304 95931
rect 163144 95869 163179 95897
rect 163207 95869 163241 95897
rect 163269 95869 163304 95897
rect 163144 95835 163304 95869
rect 163144 95807 163179 95835
rect 163207 95807 163241 95835
rect 163269 95807 163304 95835
rect 163144 95773 163304 95807
rect 163144 95745 163179 95773
rect 163207 95745 163241 95773
rect 163269 95745 163304 95773
rect 163144 95728 163304 95745
rect 178504 95959 178664 95976
rect 178504 95931 178539 95959
rect 178567 95931 178601 95959
rect 178629 95931 178664 95959
rect 178504 95897 178664 95931
rect 178504 95869 178539 95897
rect 178567 95869 178601 95897
rect 178629 95869 178664 95897
rect 178504 95835 178664 95869
rect 178504 95807 178539 95835
rect 178567 95807 178601 95835
rect 178629 95807 178664 95835
rect 178504 95773 178664 95807
rect 178504 95745 178539 95773
rect 178567 95745 178601 95773
rect 178629 95745 178664 95773
rect 178504 95728 178664 95745
rect 193864 95959 194024 95976
rect 193864 95931 193899 95959
rect 193927 95931 193961 95959
rect 193989 95931 194024 95959
rect 193864 95897 194024 95931
rect 193864 95869 193899 95897
rect 193927 95869 193961 95897
rect 193989 95869 194024 95897
rect 193864 95835 194024 95869
rect 193864 95807 193899 95835
rect 193927 95807 193961 95835
rect 193989 95807 194024 95835
rect 193864 95773 194024 95807
rect 193864 95745 193899 95773
rect 193927 95745 193961 95773
rect 193989 95745 194024 95773
rect 193864 95728 194024 95745
rect 209224 95959 209384 95976
rect 209224 95931 209259 95959
rect 209287 95931 209321 95959
rect 209349 95931 209384 95959
rect 209224 95897 209384 95931
rect 209224 95869 209259 95897
rect 209287 95869 209321 95897
rect 209349 95869 209384 95897
rect 209224 95835 209384 95869
rect 209224 95807 209259 95835
rect 209287 95807 209321 95835
rect 209349 95807 209384 95835
rect 209224 95773 209384 95807
rect 209224 95745 209259 95773
rect 209287 95745 209321 95773
rect 209349 95745 209384 95773
rect 209224 95728 209384 95745
rect 224584 95959 224744 95976
rect 224584 95931 224619 95959
rect 224647 95931 224681 95959
rect 224709 95931 224744 95959
rect 224584 95897 224744 95931
rect 224584 95869 224619 95897
rect 224647 95869 224681 95897
rect 224709 95869 224744 95897
rect 224584 95835 224744 95869
rect 224584 95807 224619 95835
rect 224647 95807 224681 95835
rect 224709 95807 224744 95835
rect 224584 95773 224744 95807
rect 224584 95745 224619 95773
rect 224647 95745 224681 95773
rect 224709 95745 224744 95773
rect 224584 95728 224744 95745
rect 239944 95959 240104 95976
rect 239944 95931 239979 95959
rect 240007 95931 240041 95959
rect 240069 95931 240104 95959
rect 239944 95897 240104 95931
rect 239944 95869 239979 95897
rect 240007 95869 240041 95897
rect 240069 95869 240104 95897
rect 239944 95835 240104 95869
rect 239944 95807 239979 95835
rect 240007 95807 240041 95835
rect 240069 95807 240104 95835
rect 239944 95773 240104 95807
rect 239944 95745 239979 95773
rect 240007 95745 240041 95773
rect 240069 95745 240104 95773
rect 239944 95728 240104 95745
rect 32584 92959 32744 92976
rect 32584 92931 32619 92959
rect 32647 92931 32681 92959
rect 32709 92931 32744 92959
rect 32584 92897 32744 92931
rect 32584 92869 32619 92897
rect 32647 92869 32681 92897
rect 32709 92869 32744 92897
rect 32584 92835 32744 92869
rect 32584 92807 32619 92835
rect 32647 92807 32681 92835
rect 32709 92807 32744 92835
rect 32584 92773 32744 92807
rect 32584 92745 32619 92773
rect 32647 92745 32681 92773
rect 32709 92745 32744 92773
rect 32584 92728 32744 92745
rect 47944 92959 48104 92976
rect 47944 92931 47979 92959
rect 48007 92931 48041 92959
rect 48069 92931 48104 92959
rect 47944 92897 48104 92931
rect 47944 92869 47979 92897
rect 48007 92869 48041 92897
rect 48069 92869 48104 92897
rect 47944 92835 48104 92869
rect 47944 92807 47979 92835
rect 48007 92807 48041 92835
rect 48069 92807 48104 92835
rect 47944 92773 48104 92807
rect 47944 92745 47979 92773
rect 48007 92745 48041 92773
rect 48069 92745 48104 92773
rect 47944 92728 48104 92745
rect 63304 92959 63464 92976
rect 63304 92931 63339 92959
rect 63367 92931 63401 92959
rect 63429 92931 63464 92959
rect 63304 92897 63464 92931
rect 63304 92869 63339 92897
rect 63367 92869 63401 92897
rect 63429 92869 63464 92897
rect 63304 92835 63464 92869
rect 63304 92807 63339 92835
rect 63367 92807 63401 92835
rect 63429 92807 63464 92835
rect 63304 92773 63464 92807
rect 63304 92745 63339 92773
rect 63367 92745 63401 92773
rect 63429 92745 63464 92773
rect 63304 92728 63464 92745
rect 78664 92959 78824 92976
rect 78664 92931 78699 92959
rect 78727 92931 78761 92959
rect 78789 92931 78824 92959
rect 78664 92897 78824 92931
rect 78664 92869 78699 92897
rect 78727 92869 78761 92897
rect 78789 92869 78824 92897
rect 78664 92835 78824 92869
rect 78664 92807 78699 92835
rect 78727 92807 78761 92835
rect 78789 92807 78824 92835
rect 78664 92773 78824 92807
rect 78664 92745 78699 92773
rect 78727 92745 78761 92773
rect 78789 92745 78824 92773
rect 78664 92728 78824 92745
rect 94024 92959 94184 92976
rect 94024 92931 94059 92959
rect 94087 92931 94121 92959
rect 94149 92931 94184 92959
rect 94024 92897 94184 92931
rect 94024 92869 94059 92897
rect 94087 92869 94121 92897
rect 94149 92869 94184 92897
rect 94024 92835 94184 92869
rect 94024 92807 94059 92835
rect 94087 92807 94121 92835
rect 94149 92807 94184 92835
rect 94024 92773 94184 92807
rect 94024 92745 94059 92773
rect 94087 92745 94121 92773
rect 94149 92745 94184 92773
rect 94024 92728 94184 92745
rect 109384 92959 109544 92976
rect 109384 92931 109419 92959
rect 109447 92931 109481 92959
rect 109509 92931 109544 92959
rect 109384 92897 109544 92931
rect 109384 92869 109419 92897
rect 109447 92869 109481 92897
rect 109509 92869 109544 92897
rect 109384 92835 109544 92869
rect 109384 92807 109419 92835
rect 109447 92807 109481 92835
rect 109509 92807 109544 92835
rect 109384 92773 109544 92807
rect 109384 92745 109419 92773
rect 109447 92745 109481 92773
rect 109509 92745 109544 92773
rect 109384 92728 109544 92745
rect 124744 92959 124904 92976
rect 124744 92931 124779 92959
rect 124807 92931 124841 92959
rect 124869 92931 124904 92959
rect 124744 92897 124904 92931
rect 124744 92869 124779 92897
rect 124807 92869 124841 92897
rect 124869 92869 124904 92897
rect 124744 92835 124904 92869
rect 124744 92807 124779 92835
rect 124807 92807 124841 92835
rect 124869 92807 124904 92835
rect 124744 92773 124904 92807
rect 124744 92745 124779 92773
rect 124807 92745 124841 92773
rect 124869 92745 124904 92773
rect 124744 92728 124904 92745
rect 140104 92959 140264 92976
rect 140104 92931 140139 92959
rect 140167 92931 140201 92959
rect 140229 92931 140264 92959
rect 140104 92897 140264 92931
rect 140104 92869 140139 92897
rect 140167 92869 140201 92897
rect 140229 92869 140264 92897
rect 140104 92835 140264 92869
rect 140104 92807 140139 92835
rect 140167 92807 140201 92835
rect 140229 92807 140264 92835
rect 140104 92773 140264 92807
rect 140104 92745 140139 92773
rect 140167 92745 140201 92773
rect 140229 92745 140264 92773
rect 140104 92728 140264 92745
rect 155464 92959 155624 92976
rect 155464 92931 155499 92959
rect 155527 92931 155561 92959
rect 155589 92931 155624 92959
rect 155464 92897 155624 92931
rect 155464 92869 155499 92897
rect 155527 92869 155561 92897
rect 155589 92869 155624 92897
rect 155464 92835 155624 92869
rect 155464 92807 155499 92835
rect 155527 92807 155561 92835
rect 155589 92807 155624 92835
rect 155464 92773 155624 92807
rect 155464 92745 155499 92773
rect 155527 92745 155561 92773
rect 155589 92745 155624 92773
rect 155464 92728 155624 92745
rect 170824 92959 170984 92976
rect 170824 92931 170859 92959
rect 170887 92931 170921 92959
rect 170949 92931 170984 92959
rect 170824 92897 170984 92931
rect 170824 92869 170859 92897
rect 170887 92869 170921 92897
rect 170949 92869 170984 92897
rect 170824 92835 170984 92869
rect 170824 92807 170859 92835
rect 170887 92807 170921 92835
rect 170949 92807 170984 92835
rect 170824 92773 170984 92807
rect 170824 92745 170859 92773
rect 170887 92745 170921 92773
rect 170949 92745 170984 92773
rect 170824 92728 170984 92745
rect 186184 92959 186344 92976
rect 186184 92931 186219 92959
rect 186247 92931 186281 92959
rect 186309 92931 186344 92959
rect 186184 92897 186344 92931
rect 186184 92869 186219 92897
rect 186247 92869 186281 92897
rect 186309 92869 186344 92897
rect 186184 92835 186344 92869
rect 186184 92807 186219 92835
rect 186247 92807 186281 92835
rect 186309 92807 186344 92835
rect 186184 92773 186344 92807
rect 186184 92745 186219 92773
rect 186247 92745 186281 92773
rect 186309 92745 186344 92773
rect 186184 92728 186344 92745
rect 201544 92959 201704 92976
rect 201544 92931 201579 92959
rect 201607 92931 201641 92959
rect 201669 92931 201704 92959
rect 201544 92897 201704 92931
rect 201544 92869 201579 92897
rect 201607 92869 201641 92897
rect 201669 92869 201704 92897
rect 201544 92835 201704 92869
rect 201544 92807 201579 92835
rect 201607 92807 201641 92835
rect 201669 92807 201704 92835
rect 201544 92773 201704 92807
rect 201544 92745 201579 92773
rect 201607 92745 201641 92773
rect 201669 92745 201704 92773
rect 201544 92728 201704 92745
rect 216904 92959 217064 92976
rect 216904 92931 216939 92959
rect 216967 92931 217001 92959
rect 217029 92931 217064 92959
rect 216904 92897 217064 92931
rect 216904 92869 216939 92897
rect 216967 92869 217001 92897
rect 217029 92869 217064 92897
rect 216904 92835 217064 92869
rect 216904 92807 216939 92835
rect 216967 92807 217001 92835
rect 217029 92807 217064 92835
rect 216904 92773 217064 92807
rect 216904 92745 216939 92773
rect 216967 92745 217001 92773
rect 217029 92745 217064 92773
rect 216904 92728 217064 92745
rect 232264 92959 232424 92976
rect 232264 92931 232299 92959
rect 232327 92931 232361 92959
rect 232389 92931 232424 92959
rect 232264 92897 232424 92931
rect 232264 92869 232299 92897
rect 232327 92869 232361 92897
rect 232389 92869 232424 92897
rect 232264 92835 232424 92869
rect 232264 92807 232299 92835
rect 232327 92807 232361 92835
rect 232389 92807 232424 92835
rect 232264 92773 232424 92807
rect 232264 92745 232299 92773
rect 232327 92745 232361 92773
rect 232389 92745 232424 92773
rect 232264 92728 232424 92745
rect 247624 92959 247784 92976
rect 247624 92931 247659 92959
rect 247687 92931 247721 92959
rect 247749 92931 247784 92959
rect 247624 92897 247784 92931
rect 247624 92869 247659 92897
rect 247687 92869 247721 92897
rect 247749 92869 247784 92897
rect 247624 92835 247784 92869
rect 247624 92807 247659 92835
rect 247687 92807 247721 92835
rect 247749 92807 247784 92835
rect 247624 92773 247784 92807
rect 247624 92745 247659 92773
rect 247687 92745 247721 92773
rect 247749 92745 247784 92773
rect 247624 92728 247784 92745
rect 254529 92959 254839 101745
rect 254529 92931 254577 92959
rect 254605 92931 254639 92959
rect 254667 92931 254701 92959
rect 254729 92931 254763 92959
rect 254791 92931 254839 92959
rect 254529 92897 254839 92931
rect 254529 92869 254577 92897
rect 254605 92869 254639 92897
rect 254667 92869 254701 92897
rect 254729 92869 254763 92897
rect 254791 92869 254839 92897
rect 254529 92835 254839 92869
rect 254529 92807 254577 92835
rect 254605 92807 254639 92835
rect 254667 92807 254701 92835
rect 254729 92807 254763 92835
rect 254791 92807 254839 92835
rect 254529 92773 254839 92807
rect 254529 92745 254577 92773
rect 254605 92745 254639 92773
rect 254667 92745 254701 92773
rect 254729 92745 254763 92773
rect 254791 92745 254839 92773
rect 31389 86931 31437 86959
rect 31465 86931 31499 86959
rect 31527 86931 31561 86959
rect 31589 86931 31623 86959
rect 31651 86931 31699 86959
rect 31389 86897 31699 86931
rect 31389 86869 31437 86897
rect 31465 86869 31499 86897
rect 31527 86869 31561 86897
rect 31589 86869 31623 86897
rect 31651 86869 31699 86897
rect 31389 86835 31699 86869
rect 31389 86807 31437 86835
rect 31465 86807 31499 86835
rect 31527 86807 31561 86835
rect 31589 86807 31623 86835
rect 31651 86807 31699 86835
rect 31389 86773 31699 86807
rect 31389 86745 31437 86773
rect 31465 86745 31499 86773
rect 31527 86745 31561 86773
rect 31589 86745 31623 86773
rect 31651 86745 31699 86773
rect 31389 77959 31699 86745
rect 40264 86959 40424 86976
rect 40264 86931 40299 86959
rect 40327 86931 40361 86959
rect 40389 86931 40424 86959
rect 40264 86897 40424 86931
rect 40264 86869 40299 86897
rect 40327 86869 40361 86897
rect 40389 86869 40424 86897
rect 40264 86835 40424 86869
rect 40264 86807 40299 86835
rect 40327 86807 40361 86835
rect 40389 86807 40424 86835
rect 40264 86773 40424 86807
rect 40264 86745 40299 86773
rect 40327 86745 40361 86773
rect 40389 86745 40424 86773
rect 40264 86728 40424 86745
rect 55624 86959 55784 86976
rect 55624 86931 55659 86959
rect 55687 86931 55721 86959
rect 55749 86931 55784 86959
rect 55624 86897 55784 86931
rect 55624 86869 55659 86897
rect 55687 86869 55721 86897
rect 55749 86869 55784 86897
rect 55624 86835 55784 86869
rect 55624 86807 55659 86835
rect 55687 86807 55721 86835
rect 55749 86807 55784 86835
rect 55624 86773 55784 86807
rect 55624 86745 55659 86773
rect 55687 86745 55721 86773
rect 55749 86745 55784 86773
rect 55624 86728 55784 86745
rect 70984 86959 71144 86976
rect 70984 86931 71019 86959
rect 71047 86931 71081 86959
rect 71109 86931 71144 86959
rect 70984 86897 71144 86931
rect 70984 86869 71019 86897
rect 71047 86869 71081 86897
rect 71109 86869 71144 86897
rect 70984 86835 71144 86869
rect 70984 86807 71019 86835
rect 71047 86807 71081 86835
rect 71109 86807 71144 86835
rect 70984 86773 71144 86807
rect 70984 86745 71019 86773
rect 71047 86745 71081 86773
rect 71109 86745 71144 86773
rect 70984 86728 71144 86745
rect 86344 86959 86504 86976
rect 86344 86931 86379 86959
rect 86407 86931 86441 86959
rect 86469 86931 86504 86959
rect 86344 86897 86504 86931
rect 86344 86869 86379 86897
rect 86407 86869 86441 86897
rect 86469 86869 86504 86897
rect 86344 86835 86504 86869
rect 86344 86807 86379 86835
rect 86407 86807 86441 86835
rect 86469 86807 86504 86835
rect 86344 86773 86504 86807
rect 86344 86745 86379 86773
rect 86407 86745 86441 86773
rect 86469 86745 86504 86773
rect 86344 86728 86504 86745
rect 101704 86959 101864 86976
rect 101704 86931 101739 86959
rect 101767 86931 101801 86959
rect 101829 86931 101864 86959
rect 101704 86897 101864 86931
rect 101704 86869 101739 86897
rect 101767 86869 101801 86897
rect 101829 86869 101864 86897
rect 101704 86835 101864 86869
rect 101704 86807 101739 86835
rect 101767 86807 101801 86835
rect 101829 86807 101864 86835
rect 101704 86773 101864 86807
rect 101704 86745 101739 86773
rect 101767 86745 101801 86773
rect 101829 86745 101864 86773
rect 101704 86728 101864 86745
rect 117064 86959 117224 86976
rect 117064 86931 117099 86959
rect 117127 86931 117161 86959
rect 117189 86931 117224 86959
rect 117064 86897 117224 86931
rect 117064 86869 117099 86897
rect 117127 86869 117161 86897
rect 117189 86869 117224 86897
rect 117064 86835 117224 86869
rect 117064 86807 117099 86835
rect 117127 86807 117161 86835
rect 117189 86807 117224 86835
rect 117064 86773 117224 86807
rect 117064 86745 117099 86773
rect 117127 86745 117161 86773
rect 117189 86745 117224 86773
rect 117064 86728 117224 86745
rect 132424 86959 132584 86976
rect 132424 86931 132459 86959
rect 132487 86931 132521 86959
rect 132549 86931 132584 86959
rect 132424 86897 132584 86931
rect 132424 86869 132459 86897
rect 132487 86869 132521 86897
rect 132549 86869 132584 86897
rect 132424 86835 132584 86869
rect 132424 86807 132459 86835
rect 132487 86807 132521 86835
rect 132549 86807 132584 86835
rect 132424 86773 132584 86807
rect 132424 86745 132459 86773
rect 132487 86745 132521 86773
rect 132549 86745 132584 86773
rect 132424 86728 132584 86745
rect 147784 86959 147944 86976
rect 147784 86931 147819 86959
rect 147847 86931 147881 86959
rect 147909 86931 147944 86959
rect 147784 86897 147944 86931
rect 147784 86869 147819 86897
rect 147847 86869 147881 86897
rect 147909 86869 147944 86897
rect 147784 86835 147944 86869
rect 147784 86807 147819 86835
rect 147847 86807 147881 86835
rect 147909 86807 147944 86835
rect 147784 86773 147944 86807
rect 147784 86745 147819 86773
rect 147847 86745 147881 86773
rect 147909 86745 147944 86773
rect 147784 86728 147944 86745
rect 163144 86959 163304 86976
rect 163144 86931 163179 86959
rect 163207 86931 163241 86959
rect 163269 86931 163304 86959
rect 163144 86897 163304 86931
rect 163144 86869 163179 86897
rect 163207 86869 163241 86897
rect 163269 86869 163304 86897
rect 163144 86835 163304 86869
rect 163144 86807 163179 86835
rect 163207 86807 163241 86835
rect 163269 86807 163304 86835
rect 163144 86773 163304 86807
rect 163144 86745 163179 86773
rect 163207 86745 163241 86773
rect 163269 86745 163304 86773
rect 163144 86728 163304 86745
rect 178504 86959 178664 86976
rect 178504 86931 178539 86959
rect 178567 86931 178601 86959
rect 178629 86931 178664 86959
rect 178504 86897 178664 86931
rect 178504 86869 178539 86897
rect 178567 86869 178601 86897
rect 178629 86869 178664 86897
rect 178504 86835 178664 86869
rect 178504 86807 178539 86835
rect 178567 86807 178601 86835
rect 178629 86807 178664 86835
rect 178504 86773 178664 86807
rect 178504 86745 178539 86773
rect 178567 86745 178601 86773
rect 178629 86745 178664 86773
rect 178504 86728 178664 86745
rect 193864 86959 194024 86976
rect 193864 86931 193899 86959
rect 193927 86931 193961 86959
rect 193989 86931 194024 86959
rect 193864 86897 194024 86931
rect 193864 86869 193899 86897
rect 193927 86869 193961 86897
rect 193989 86869 194024 86897
rect 193864 86835 194024 86869
rect 193864 86807 193899 86835
rect 193927 86807 193961 86835
rect 193989 86807 194024 86835
rect 193864 86773 194024 86807
rect 193864 86745 193899 86773
rect 193927 86745 193961 86773
rect 193989 86745 194024 86773
rect 193864 86728 194024 86745
rect 209224 86959 209384 86976
rect 209224 86931 209259 86959
rect 209287 86931 209321 86959
rect 209349 86931 209384 86959
rect 209224 86897 209384 86931
rect 209224 86869 209259 86897
rect 209287 86869 209321 86897
rect 209349 86869 209384 86897
rect 209224 86835 209384 86869
rect 209224 86807 209259 86835
rect 209287 86807 209321 86835
rect 209349 86807 209384 86835
rect 209224 86773 209384 86807
rect 209224 86745 209259 86773
rect 209287 86745 209321 86773
rect 209349 86745 209384 86773
rect 209224 86728 209384 86745
rect 224584 86959 224744 86976
rect 224584 86931 224619 86959
rect 224647 86931 224681 86959
rect 224709 86931 224744 86959
rect 224584 86897 224744 86931
rect 224584 86869 224619 86897
rect 224647 86869 224681 86897
rect 224709 86869 224744 86897
rect 224584 86835 224744 86869
rect 224584 86807 224619 86835
rect 224647 86807 224681 86835
rect 224709 86807 224744 86835
rect 224584 86773 224744 86807
rect 224584 86745 224619 86773
rect 224647 86745 224681 86773
rect 224709 86745 224744 86773
rect 224584 86728 224744 86745
rect 239944 86959 240104 86976
rect 239944 86931 239979 86959
rect 240007 86931 240041 86959
rect 240069 86931 240104 86959
rect 239944 86897 240104 86931
rect 239944 86869 239979 86897
rect 240007 86869 240041 86897
rect 240069 86869 240104 86897
rect 239944 86835 240104 86869
rect 239944 86807 239979 86835
rect 240007 86807 240041 86835
rect 240069 86807 240104 86835
rect 239944 86773 240104 86807
rect 239944 86745 239979 86773
rect 240007 86745 240041 86773
rect 240069 86745 240104 86773
rect 239944 86728 240104 86745
rect 32584 83959 32744 83976
rect 32584 83931 32619 83959
rect 32647 83931 32681 83959
rect 32709 83931 32744 83959
rect 32584 83897 32744 83931
rect 32584 83869 32619 83897
rect 32647 83869 32681 83897
rect 32709 83869 32744 83897
rect 32584 83835 32744 83869
rect 32584 83807 32619 83835
rect 32647 83807 32681 83835
rect 32709 83807 32744 83835
rect 32584 83773 32744 83807
rect 32584 83745 32619 83773
rect 32647 83745 32681 83773
rect 32709 83745 32744 83773
rect 32584 83728 32744 83745
rect 47944 83959 48104 83976
rect 47944 83931 47979 83959
rect 48007 83931 48041 83959
rect 48069 83931 48104 83959
rect 47944 83897 48104 83931
rect 47944 83869 47979 83897
rect 48007 83869 48041 83897
rect 48069 83869 48104 83897
rect 47944 83835 48104 83869
rect 47944 83807 47979 83835
rect 48007 83807 48041 83835
rect 48069 83807 48104 83835
rect 47944 83773 48104 83807
rect 47944 83745 47979 83773
rect 48007 83745 48041 83773
rect 48069 83745 48104 83773
rect 47944 83728 48104 83745
rect 63304 83959 63464 83976
rect 63304 83931 63339 83959
rect 63367 83931 63401 83959
rect 63429 83931 63464 83959
rect 63304 83897 63464 83931
rect 63304 83869 63339 83897
rect 63367 83869 63401 83897
rect 63429 83869 63464 83897
rect 63304 83835 63464 83869
rect 63304 83807 63339 83835
rect 63367 83807 63401 83835
rect 63429 83807 63464 83835
rect 63304 83773 63464 83807
rect 63304 83745 63339 83773
rect 63367 83745 63401 83773
rect 63429 83745 63464 83773
rect 63304 83728 63464 83745
rect 78664 83959 78824 83976
rect 78664 83931 78699 83959
rect 78727 83931 78761 83959
rect 78789 83931 78824 83959
rect 78664 83897 78824 83931
rect 78664 83869 78699 83897
rect 78727 83869 78761 83897
rect 78789 83869 78824 83897
rect 78664 83835 78824 83869
rect 78664 83807 78699 83835
rect 78727 83807 78761 83835
rect 78789 83807 78824 83835
rect 78664 83773 78824 83807
rect 78664 83745 78699 83773
rect 78727 83745 78761 83773
rect 78789 83745 78824 83773
rect 78664 83728 78824 83745
rect 94024 83959 94184 83976
rect 94024 83931 94059 83959
rect 94087 83931 94121 83959
rect 94149 83931 94184 83959
rect 94024 83897 94184 83931
rect 94024 83869 94059 83897
rect 94087 83869 94121 83897
rect 94149 83869 94184 83897
rect 94024 83835 94184 83869
rect 94024 83807 94059 83835
rect 94087 83807 94121 83835
rect 94149 83807 94184 83835
rect 94024 83773 94184 83807
rect 94024 83745 94059 83773
rect 94087 83745 94121 83773
rect 94149 83745 94184 83773
rect 94024 83728 94184 83745
rect 109384 83959 109544 83976
rect 109384 83931 109419 83959
rect 109447 83931 109481 83959
rect 109509 83931 109544 83959
rect 109384 83897 109544 83931
rect 109384 83869 109419 83897
rect 109447 83869 109481 83897
rect 109509 83869 109544 83897
rect 109384 83835 109544 83869
rect 109384 83807 109419 83835
rect 109447 83807 109481 83835
rect 109509 83807 109544 83835
rect 109384 83773 109544 83807
rect 109384 83745 109419 83773
rect 109447 83745 109481 83773
rect 109509 83745 109544 83773
rect 109384 83728 109544 83745
rect 124744 83959 124904 83976
rect 124744 83931 124779 83959
rect 124807 83931 124841 83959
rect 124869 83931 124904 83959
rect 124744 83897 124904 83931
rect 124744 83869 124779 83897
rect 124807 83869 124841 83897
rect 124869 83869 124904 83897
rect 124744 83835 124904 83869
rect 124744 83807 124779 83835
rect 124807 83807 124841 83835
rect 124869 83807 124904 83835
rect 124744 83773 124904 83807
rect 124744 83745 124779 83773
rect 124807 83745 124841 83773
rect 124869 83745 124904 83773
rect 124744 83728 124904 83745
rect 140104 83959 140264 83976
rect 140104 83931 140139 83959
rect 140167 83931 140201 83959
rect 140229 83931 140264 83959
rect 140104 83897 140264 83931
rect 140104 83869 140139 83897
rect 140167 83869 140201 83897
rect 140229 83869 140264 83897
rect 140104 83835 140264 83869
rect 140104 83807 140139 83835
rect 140167 83807 140201 83835
rect 140229 83807 140264 83835
rect 140104 83773 140264 83807
rect 140104 83745 140139 83773
rect 140167 83745 140201 83773
rect 140229 83745 140264 83773
rect 140104 83728 140264 83745
rect 155464 83959 155624 83976
rect 155464 83931 155499 83959
rect 155527 83931 155561 83959
rect 155589 83931 155624 83959
rect 155464 83897 155624 83931
rect 155464 83869 155499 83897
rect 155527 83869 155561 83897
rect 155589 83869 155624 83897
rect 155464 83835 155624 83869
rect 155464 83807 155499 83835
rect 155527 83807 155561 83835
rect 155589 83807 155624 83835
rect 155464 83773 155624 83807
rect 155464 83745 155499 83773
rect 155527 83745 155561 83773
rect 155589 83745 155624 83773
rect 155464 83728 155624 83745
rect 170824 83959 170984 83976
rect 170824 83931 170859 83959
rect 170887 83931 170921 83959
rect 170949 83931 170984 83959
rect 170824 83897 170984 83931
rect 170824 83869 170859 83897
rect 170887 83869 170921 83897
rect 170949 83869 170984 83897
rect 170824 83835 170984 83869
rect 170824 83807 170859 83835
rect 170887 83807 170921 83835
rect 170949 83807 170984 83835
rect 170824 83773 170984 83807
rect 170824 83745 170859 83773
rect 170887 83745 170921 83773
rect 170949 83745 170984 83773
rect 170824 83728 170984 83745
rect 186184 83959 186344 83976
rect 186184 83931 186219 83959
rect 186247 83931 186281 83959
rect 186309 83931 186344 83959
rect 186184 83897 186344 83931
rect 186184 83869 186219 83897
rect 186247 83869 186281 83897
rect 186309 83869 186344 83897
rect 186184 83835 186344 83869
rect 186184 83807 186219 83835
rect 186247 83807 186281 83835
rect 186309 83807 186344 83835
rect 186184 83773 186344 83807
rect 186184 83745 186219 83773
rect 186247 83745 186281 83773
rect 186309 83745 186344 83773
rect 186184 83728 186344 83745
rect 201544 83959 201704 83976
rect 201544 83931 201579 83959
rect 201607 83931 201641 83959
rect 201669 83931 201704 83959
rect 201544 83897 201704 83931
rect 201544 83869 201579 83897
rect 201607 83869 201641 83897
rect 201669 83869 201704 83897
rect 201544 83835 201704 83869
rect 201544 83807 201579 83835
rect 201607 83807 201641 83835
rect 201669 83807 201704 83835
rect 201544 83773 201704 83807
rect 201544 83745 201579 83773
rect 201607 83745 201641 83773
rect 201669 83745 201704 83773
rect 201544 83728 201704 83745
rect 216904 83959 217064 83976
rect 216904 83931 216939 83959
rect 216967 83931 217001 83959
rect 217029 83931 217064 83959
rect 216904 83897 217064 83931
rect 216904 83869 216939 83897
rect 216967 83869 217001 83897
rect 217029 83869 217064 83897
rect 216904 83835 217064 83869
rect 216904 83807 216939 83835
rect 216967 83807 217001 83835
rect 217029 83807 217064 83835
rect 216904 83773 217064 83807
rect 216904 83745 216939 83773
rect 216967 83745 217001 83773
rect 217029 83745 217064 83773
rect 216904 83728 217064 83745
rect 232264 83959 232424 83976
rect 232264 83931 232299 83959
rect 232327 83931 232361 83959
rect 232389 83931 232424 83959
rect 232264 83897 232424 83931
rect 232264 83869 232299 83897
rect 232327 83869 232361 83897
rect 232389 83869 232424 83897
rect 232264 83835 232424 83869
rect 232264 83807 232299 83835
rect 232327 83807 232361 83835
rect 232389 83807 232424 83835
rect 232264 83773 232424 83807
rect 232264 83745 232299 83773
rect 232327 83745 232361 83773
rect 232389 83745 232424 83773
rect 232264 83728 232424 83745
rect 247624 83959 247784 83976
rect 247624 83931 247659 83959
rect 247687 83931 247721 83959
rect 247749 83931 247784 83959
rect 247624 83897 247784 83931
rect 247624 83869 247659 83897
rect 247687 83869 247721 83897
rect 247749 83869 247784 83897
rect 247624 83835 247784 83869
rect 247624 83807 247659 83835
rect 247687 83807 247721 83835
rect 247749 83807 247784 83835
rect 247624 83773 247784 83807
rect 247624 83745 247659 83773
rect 247687 83745 247721 83773
rect 247749 83745 247784 83773
rect 247624 83728 247784 83745
rect 254529 83959 254839 92745
rect 254529 83931 254577 83959
rect 254605 83931 254639 83959
rect 254667 83931 254701 83959
rect 254729 83931 254763 83959
rect 254791 83931 254839 83959
rect 254529 83897 254839 83931
rect 254529 83869 254577 83897
rect 254605 83869 254639 83897
rect 254667 83869 254701 83897
rect 254729 83869 254763 83897
rect 254791 83869 254839 83897
rect 254529 83835 254839 83869
rect 254529 83807 254577 83835
rect 254605 83807 254639 83835
rect 254667 83807 254701 83835
rect 254729 83807 254763 83835
rect 254791 83807 254839 83835
rect 254529 83773 254839 83807
rect 254529 83745 254577 83773
rect 254605 83745 254639 83773
rect 254667 83745 254701 83773
rect 254729 83745 254763 83773
rect 254791 83745 254839 83773
rect 31389 77931 31437 77959
rect 31465 77931 31499 77959
rect 31527 77931 31561 77959
rect 31589 77931 31623 77959
rect 31651 77931 31699 77959
rect 31389 77897 31699 77931
rect 31389 77869 31437 77897
rect 31465 77869 31499 77897
rect 31527 77869 31561 77897
rect 31589 77869 31623 77897
rect 31651 77869 31699 77897
rect 31389 77835 31699 77869
rect 31389 77807 31437 77835
rect 31465 77807 31499 77835
rect 31527 77807 31561 77835
rect 31589 77807 31623 77835
rect 31651 77807 31699 77835
rect 31389 77773 31699 77807
rect 31389 77745 31437 77773
rect 31465 77745 31499 77773
rect 31527 77745 31561 77773
rect 31589 77745 31623 77773
rect 31651 77745 31699 77773
rect 31389 68959 31699 77745
rect 40264 77959 40424 77976
rect 40264 77931 40299 77959
rect 40327 77931 40361 77959
rect 40389 77931 40424 77959
rect 40264 77897 40424 77931
rect 40264 77869 40299 77897
rect 40327 77869 40361 77897
rect 40389 77869 40424 77897
rect 40264 77835 40424 77869
rect 40264 77807 40299 77835
rect 40327 77807 40361 77835
rect 40389 77807 40424 77835
rect 40264 77773 40424 77807
rect 40264 77745 40299 77773
rect 40327 77745 40361 77773
rect 40389 77745 40424 77773
rect 40264 77728 40424 77745
rect 55624 77959 55784 77976
rect 55624 77931 55659 77959
rect 55687 77931 55721 77959
rect 55749 77931 55784 77959
rect 55624 77897 55784 77931
rect 55624 77869 55659 77897
rect 55687 77869 55721 77897
rect 55749 77869 55784 77897
rect 55624 77835 55784 77869
rect 55624 77807 55659 77835
rect 55687 77807 55721 77835
rect 55749 77807 55784 77835
rect 55624 77773 55784 77807
rect 55624 77745 55659 77773
rect 55687 77745 55721 77773
rect 55749 77745 55784 77773
rect 55624 77728 55784 77745
rect 70984 77959 71144 77976
rect 70984 77931 71019 77959
rect 71047 77931 71081 77959
rect 71109 77931 71144 77959
rect 70984 77897 71144 77931
rect 70984 77869 71019 77897
rect 71047 77869 71081 77897
rect 71109 77869 71144 77897
rect 70984 77835 71144 77869
rect 70984 77807 71019 77835
rect 71047 77807 71081 77835
rect 71109 77807 71144 77835
rect 70984 77773 71144 77807
rect 70984 77745 71019 77773
rect 71047 77745 71081 77773
rect 71109 77745 71144 77773
rect 70984 77728 71144 77745
rect 86344 77959 86504 77976
rect 86344 77931 86379 77959
rect 86407 77931 86441 77959
rect 86469 77931 86504 77959
rect 86344 77897 86504 77931
rect 86344 77869 86379 77897
rect 86407 77869 86441 77897
rect 86469 77869 86504 77897
rect 86344 77835 86504 77869
rect 86344 77807 86379 77835
rect 86407 77807 86441 77835
rect 86469 77807 86504 77835
rect 86344 77773 86504 77807
rect 86344 77745 86379 77773
rect 86407 77745 86441 77773
rect 86469 77745 86504 77773
rect 86344 77728 86504 77745
rect 101704 77959 101864 77976
rect 101704 77931 101739 77959
rect 101767 77931 101801 77959
rect 101829 77931 101864 77959
rect 101704 77897 101864 77931
rect 101704 77869 101739 77897
rect 101767 77869 101801 77897
rect 101829 77869 101864 77897
rect 101704 77835 101864 77869
rect 101704 77807 101739 77835
rect 101767 77807 101801 77835
rect 101829 77807 101864 77835
rect 101704 77773 101864 77807
rect 101704 77745 101739 77773
rect 101767 77745 101801 77773
rect 101829 77745 101864 77773
rect 101704 77728 101864 77745
rect 117064 77959 117224 77976
rect 117064 77931 117099 77959
rect 117127 77931 117161 77959
rect 117189 77931 117224 77959
rect 117064 77897 117224 77931
rect 117064 77869 117099 77897
rect 117127 77869 117161 77897
rect 117189 77869 117224 77897
rect 117064 77835 117224 77869
rect 117064 77807 117099 77835
rect 117127 77807 117161 77835
rect 117189 77807 117224 77835
rect 117064 77773 117224 77807
rect 117064 77745 117099 77773
rect 117127 77745 117161 77773
rect 117189 77745 117224 77773
rect 117064 77728 117224 77745
rect 132424 77959 132584 77976
rect 132424 77931 132459 77959
rect 132487 77931 132521 77959
rect 132549 77931 132584 77959
rect 132424 77897 132584 77931
rect 132424 77869 132459 77897
rect 132487 77869 132521 77897
rect 132549 77869 132584 77897
rect 132424 77835 132584 77869
rect 132424 77807 132459 77835
rect 132487 77807 132521 77835
rect 132549 77807 132584 77835
rect 132424 77773 132584 77807
rect 132424 77745 132459 77773
rect 132487 77745 132521 77773
rect 132549 77745 132584 77773
rect 132424 77728 132584 77745
rect 147784 77959 147944 77976
rect 147784 77931 147819 77959
rect 147847 77931 147881 77959
rect 147909 77931 147944 77959
rect 147784 77897 147944 77931
rect 147784 77869 147819 77897
rect 147847 77869 147881 77897
rect 147909 77869 147944 77897
rect 147784 77835 147944 77869
rect 147784 77807 147819 77835
rect 147847 77807 147881 77835
rect 147909 77807 147944 77835
rect 147784 77773 147944 77807
rect 147784 77745 147819 77773
rect 147847 77745 147881 77773
rect 147909 77745 147944 77773
rect 147784 77728 147944 77745
rect 163144 77959 163304 77976
rect 163144 77931 163179 77959
rect 163207 77931 163241 77959
rect 163269 77931 163304 77959
rect 163144 77897 163304 77931
rect 163144 77869 163179 77897
rect 163207 77869 163241 77897
rect 163269 77869 163304 77897
rect 163144 77835 163304 77869
rect 163144 77807 163179 77835
rect 163207 77807 163241 77835
rect 163269 77807 163304 77835
rect 163144 77773 163304 77807
rect 163144 77745 163179 77773
rect 163207 77745 163241 77773
rect 163269 77745 163304 77773
rect 163144 77728 163304 77745
rect 178504 77959 178664 77976
rect 178504 77931 178539 77959
rect 178567 77931 178601 77959
rect 178629 77931 178664 77959
rect 178504 77897 178664 77931
rect 178504 77869 178539 77897
rect 178567 77869 178601 77897
rect 178629 77869 178664 77897
rect 178504 77835 178664 77869
rect 178504 77807 178539 77835
rect 178567 77807 178601 77835
rect 178629 77807 178664 77835
rect 178504 77773 178664 77807
rect 178504 77745 178539 77773
rect 178567 77745 178601 77773
rect 178629 77745 178664 77773
rect 178504 77728 178664 77745
rect 193864 77959 194024 77976
rect 193864 77931 193899 77959
rect 193927 77931 193961 77959
rect 193989 77931 194024 77959
rect 193864 77897 194024 77931
rect 193864 77869 193899 77897
rect 193927 77869 193961 77897
rect 193989 77869 194024 77897
rect 193864 77835 194024 77869
rect 193864 77807 193899 77835
rect 193927 77807 193961 77835
rect 193989 77807 194024 77835
rect 193864 77773 194024 77807
rect 193864 77745 193899 77773
rect 193927 77745 193961 77773
rect 193989 77745 194024 77773
rect 193864 77728 194024 77745
rect 209224 77959 209384 77976
rect 209224 77931 209259 77959
rect 209287 77931 209321 77959
rect 209349 77931 209384 77959
rect 209224 77897 209384 77931
rect 209224 77869 209259 77897
rect 209287 77869 209321 77897
rect 209349 77869 209384 77897
rect 209224 77835 209384 77869
rect 209224 77807 209259 77835
rect 209287 77807 209321 77835
rect 209349 77807 209384 77835
rect 209224 77773 209384 77807
rect 209224 77745 209259 77773
rect 209287 77745 209321 77773
rect 209349 77745 209384 77773
rect 209224 77728 209384 77745
rect 224584 77959 224744 77976
rect 224584 77931 224619 77959
rect 224647 77931 224681 77959
rect 224709 77931 224744 77959
rect 224584 77897 224744 77931
rect 224584 77869 224619 77897
rect 224647 77869 224681 77897
rect 224709 77869 224744 77897
rect 224584 77835 224744 77869
rect 224584 77807 224619 77835
rect 224647 77807 224681 77835
rect 224709 77807 224744 77835
rect 224584 77773 224744 77807
rect 224584 77745 224619 77773
rect 224647 77745 224681 77773
rect 224709 77745 224744 77773
rect 224584 77728 224744 77745
rect 239944 77959 240104 77976
rect 239944 77931 239979 77959
rect 240007 77931 240041 77959
rect 240069 77931 240104 77959
rect 239944 77897 240104 77931
rect 239944 77869 239979 77897
rect 240007 77869 240041 77897
rect 240069 77869 240104 77897
rect 239944 77835 240104 77869
rect 239944 77807 239979 77835
rect 240007 77807 240041 77835
rect 240069 77807 240104 77835
rect 239944 77773 240104 77807
rect 239944 77745 239979 77773
rect 240007 77745 240041 77773
rect 240069 77745 240104 77773
rect 239944 77728 240104 77745
rect 32584 74959 32744 74976
rect 32584 74931 32619 74959
rect 32647 74931 32681 74959
rect 32709 74931 32744 74959
rect 32584 74897 32744 74931
rect 32584 74869 32619 74897
rect 32647 74869 32681 74897
rect 32709 74869 32744 74897
rect 32584 74835 32744 74869
rect 32584 74807 32619 74835
rect 32647 74807 32681 74835
rect 32709 74807 32744 74835
rect 32584 74773 32744 74807
rect 32584 74745 32619 74773
rect 32647 74745 32681 74773
rect 32709 74745 32744 74773
rect 32584 74728 32744 74745
rect 47944 74959 48104 74976
rect 47944 74931 47979 74959
rect 48007 74931 48041 74959
rect 48069 74931 48104 74959
rect 47944 74897 48104 74931
rect 47944 74869 47979 74897
rect 48007 74869 48041 74897
rect 48069 74869 48104 74897
rect 47944 74835 48104 74869
rect 47944 74807 47979 74835
rect 48007 74807 48041 74835
rect 48069 74807 48104 74835
rect 47944 74773 48104 74807
rect 47944 74745 47979 74773
rect 48007 74745 48041 74773
rect 48069 74745 48104 74773
rect 47944 74728 48104 74745
rect 63304 74959 63464 74976
rect 63304 74931 63339 74959
rect 63367 74931 63401 74959
rect 63429 74931 63464 74959
rect 63304 74897 63464 74931
rect 63304 74869 63339 74897
rect 63367 74869 63401 74897
rect 63429 74869 63464 74897
rect 63304 74835 63464 74869
rect 63304 74807 63339 74835
rect 63367 74807 63401 74835
rect 63429 74807 63464 74835
rect 63304 74773 63464 74807
rect 63304 74745 63339 74773
rect 63367 74745 63401 74773
rect 63429 74745 63464 74773
rect 63304 74728 63464 74745
rect 78664 74959 78824 74976
rect 78664 74931 78699 74959
rect 78727 74931 78761 74959
rect 78789 74931 78824 74959
rect 78664 74897 78824 74931
rect 78664 74869 78699 74897
rect 78727 74869 78761 74897
rect 78789 74869 78824 74897
rect 78664 74835 78824 74869
rect 78664 74807 78699 74835
rect 78727 74807 78761 74835
rect 78789 74807 78824 74835
rect 78664 74773 78824 74807
rect 78664 74745 78699 74773
rect 78727 74745 78761 74773
rect 78789 74745 78824 74773
rect 78664 74728 78824 74745
rect 94024 74959 94184 74976
rect 94024 74931 94059 74959
rect 94087 74931 94121 74959
rect 94149 74931 94184 74959
rect 94024 74897 94184 74931
rect 94024 74869 94059 74897
rect 94087 74869 94121 74897
rect 94149 74869 94184 74897
rect 94024 74835 94184 74869
rect 94024 74807 94059 74835
rect 94087 74807 94121 74835
rect 94149 74807 94184 74835
rect 94024 74773 94184 74807
rect 94024 74745 94059 74773
rect 94087 74745 94121 74773
rect 94149 74745 94184 74773
rect 94024 74728 94184 74745
rect 109384 74959 109544 74976
rect 109384 74931 109419 74959
rect 109447 74931 109481 74959
rect 109509 74931 109544 74959
rect 109384 74897 109544 74931
rect 109384 74869 109419 74897
rect 109447 74869 109481 74897
rect 109509 74869 109544 74897
rect 109384 74835 109544 74869
rect 109384 74807 109419 74835
rect 109447 74807 109481 74835
rect 109509 74807 109544 74835
rect 109384 74773 109544 74807
rect 109384 74745 109419 74773
rect 109447 74745 109481 74773
rect 109509 74745 109544 74773
rect 109384 74728 109544 74745
rect 124744 74959 124904 74976
rect 124744 74931 124779 74959
rect 124807 74931 124841 74959
rect 124869 74931 124904 74959
rect 124744 74897 124904 74931
rect 124744 74869 124779 74897
rect 124807 74869 124841 74897
rect 124869 74869 124904 74897
rect 124744 74835 124904 74869
rect 124744 74807 124779 74835
rect 124807 74807 124841 74835
rect 124869 74807 124904 74835
rect 124744 74773 124904 74807
rect 124744 74745 124779 74773
rect 124807 74745 124841 74773
rect 124869 74745 124904 74773
rect 124744 74728 124904 74745
rect 140104 74959 140264 74976
rect 140104 74931 140139 74959
rect 140167 74931 140201 74959
rect 140229 74931 140264 74959
rect 140104 74897 140264 74931
rect 140104 74869 140139 74897
rect 140167 74869 140201 74897
rect 140229 74869 140264 74897
rect 140104 74835 140264 74869
rect 140104 74807 140139 74835
rect 140167 74807 140201 74835
rect 140229 74807 140264 74835
rect 140104 74773 140264 74807
rect 140104 74745 140139 74773
rect 140167 74745 140201 74773
rect 140229 74745 140264 74773
rect 140104 74728 140264 74745
rect 155464 74959 155624 74976
rect 155464 74931 155499 74959
rect 155527 74931 155561 74959
rect 155589 74931 155624 74959
rect 155464 74897 155624 74931
rect 155464 74869 155499 74897
rect 155527 74869 155561 74897
rect 155589 74869 155624 74897
rect 155464 74835 155624 74869
rect 155464 74807 155499 74835
rect 155527 74807 155561 74835
rect 155589 74807 155624 74835
rect 155464 74773 155624 74807
rect 155464 74745 155499 74773
rect 155527 74745 155561 74773
rect 155589 74745 155624 74773
rect 155464 74728 155624 74745
rect 170824 74959 170984 74976
rect 170824 74931 170859 74959
rect 170887 74931 170921 74959
rect 170949 74931 170984 74959
rect 170824 74897 170984 74931
rect 170824 74869 170859 74897
rect 170887 74869 170921 74897
rect 170949 74869 170984 74897
rect 170824 74835 170984 74869
rect 170824 74807 170859 74835
rect 170887 74807 170921 74835
rect 170949 74807 170984 74835
rect 170824 74773 170984 74807
rect 170824 74745 170859 74773
rect 170887 74745 170921 74773
rect 170949 74745 170984 74773
rect 170824 74728 170984 74745
rect 186184 74959 186344 74976
rect 186184 74931 186219 74959
rect 186247 74931 186281 74959
rect 186309 74931 186344 74959
rect 186184 74897 186344 74931
rect 186184 74869 186219 74897
rect 186247 74869 186281 74897
rect 186309 74869 186344 74897
rect 186184 74835 186344 74869
rect 186184 74807 186219 74835
rect 186247 74807 186281 74835
rect 186309 74807 186344 74835
rect 186184 74773 186344 74807
rect 186184 74745 186219 74773
rect 186247 74745 186281 74773
rect 186309 74745 186344 74773
rect 186184 74728 186344 74745
rect 201544 74959 201704 74976
rect 201544 74931 201579 74959
rect 201607 74931 201641 74959
rect 201669 74931 201704 74959
rect 201544 74897 201704 74931
rect 201544 74869 201579 74897
rect 201607 74869 201641 74897
rect 201669 74869 201704 74897
rect 201544 74835 201704 74869
rect 201544 74807 201579 74835
rect 201607 74807 201641 74835
rect 201669 74807 201704 74835
rect 201544 74773 201704 74807
rect 201544 74745 201579 74773
rect 201607 74745 201641 74773
rect 201669 74745 201704 74773
rect 201544 74728 201704 74745
rect 216904 74959 217064 74976
rect 216904 74931 216939 74959
rect 216967 74931 217001 74959
rect 217029 74931 217064 74959
rect 216904 74897 217064 74931
rect 216904 74869 216939 74897
rect 216967 74869 217001 74897
rect 217029 74869 217064 74897
rect 216904 74835 217064 74869
rect 216904 74807 216939 74835
rect 216967 74807 217001 74835
rect 217029 74807 217064 74835
rect 216904 74773 217064 74807
rect 216904 74745 216939 74773
rect 216967 74745 217001 74773
rect 217029 74745 217064 74773
rect 216904 74728 217064 74745
rect 232264 74959 232424 74976
rect 232264 74931 232299 74959
rect 232327 74931 232361 74959
rect 232389 74931 232424 74959
rect 232264 74897 232424 74931
rect 232264 74869 232299 74897
rect 232327 74869 232361 74897
rect 232389 74869 232424 74897
rect 232264 74835 232424 74869
rect 232264 74807 232299 74835
rect 232327 74807 232361 74835
rect 232389 74807 232424 74835
rect 232264 74773 232424 74807
rect 232264 74745 232299 74773
rect 232327 74745 232361 74773
rect 232389 74745 232424 74773
rect 232264 74728 232424 74745
rect 247624 74959 247784 74976
rect 247624 74931 247659 74959
rect 247687 74931 247721 74959
rect 247749 74931 247784 74959
rect 247624 74897 247784 74931
rect 247624 74869 247659 74897
rect 247687 74869 247721 74897
rect 247749 74869 247784 74897
rect 247624 74835 247784 74869
rect 247624 74807 247659 74835
rect 247687 74807 247721 74835
rect 247749 74807 247784 74835
rect 247624 74773 247784 74807
rect 247624 74745 247659 74773
rect 247687 74745 247721 74773
rect 247749 74745 247784 74773
rect 247624 74728 247784 74745
rect 254529 74959 254839 83745
rect 254529 74931 254577 74959
rect 254605 74931 254639 74959
rect 254667 74931 254701 74959
rect 254729 74931 254763 74959
rect 254791 74931 254839 74959
rect 254529 74897 254839 74931
rect 254529 74869 254577 74897
rect 254605 74869 254639 74897
rect 254667 74869 254701 74897
rect 254729 74869 254763 74897
rect 254791 74869 254839 74897
rect 254529 74835 254839 74869
rect 254529 74807 254577 74835
rect 254605 74807 254639 74835
rect 254667 74807 254701 74835
rect 254729 74807 254763 74835
rect 254791 74807 254839 74835
rect 254529 74773 254839 74807
rect 254529 74745 254577 74773
rect 254605 74745 254639 74773
rect 254667 74745 254701 74773
rect 254729 74745 254763 74773
rect 254791 74745 254839 74773
rect 31389 68931 31437 68959
rect 31465 68931 31499 68959
rect 31527 68931 31561 68959
rect 31589 68931 31623 68959
rect 31651 68931 31699 68959
rect 31389 68897 31699 68931
rect 31389 68869 31437 68897
rect 31465 68869 31499 68897
rect 31527 68869 31561 68897
rect 31589 68869 31623 68897
rect 31651 68869 31699 68897
rect 31389 68835 31699 68869
rect 31389 68807 31437 68835
rect 31465 68807 31499 68835
rect 31527 68807 31561 68835
rect 31589 68807 31623 68835
rect 31651 68807 31699 68835
rect 31389 68773 31699 68807
rect 31389 68745 31437 68773
rect 31465 68745 31499 68773
rect 31527 68745 31561 68773
rect 31589 68745 31623 68773
rect 31651 68745 31699 68773
rect 31389 59959 31699 68745
rect 40264 68959 40424 68976
rect 40264 68931 40299 68959
rect 40327 68931 40361 68959
rect 40389 68931 40424 68959
rect 40264 68897 40424 68931
rect 40264 68869 40299 68897
rect 40327 68869 40361 68897
rect 40389 68869 40424 68897
rect 40264 68835 40424 68869
rect 40264 68807 40299 68835
rect 40327 68807 40361 68835
rect 40389 68807 40424 68835
rect 40264 68773 40424 68807
rect 40264 68745 40299 68773
rect 40327 68745 40361 68773
rect 40389 68745 40424 68773
rect 40264 68728 40424 68745
rect 55624 68959 55784 68976
rect 55624 68931 55659 68959
rect 55687 68931 55721 68959
rect 55749 68931 55784 68959
rect 55624 68897 55784 68931
rect 55624 68869 55659 68897
rect 55687 68869 55721 68897
rect 55749 68869 55784 68897
rect 55624 68835 55784 68869
rect 55624 68807 55659 68835
rect 55687 68807 55721 68835
rect 55749 68807 55784 68835
rect 55624 68773 55784 68807
rect 55624 68745 55659 68773
rect 55687 68745 55721 68773
rect 55749 68745 55784 68773
rect 55624 68728 55784 68745
rect 70984 68959 71144 68976
rect 70984 68931 71019 68959
rect 71047 68931 71081 68959
rect 71109 68931 71144 68959
rect 70984 68897 71144 68931
rect 70984 68869 71019 68897
rect 71047 68869 71081 68897
rect 71109 68869 71144 68897
rect 70984 68835 71144 68869
rect 70984 68807 71019 68835
rect 71047 68807 71081 68835
rect 71109 68807 71144 68835
rect 70984 68773 71144 68807
rect 70984 68745 71019 68773
rect 71047 68745 71081 68773
rect 71109 68745 71144 68773
rect 70984 68728 71144 68745
rect 86344 68959 86504 68976
rect 86344 68931 86379 68959
rect 86407 68931 86441 68959
rect 86469 68931 86504 68959
rect 86344 68897 86504 68931
rect 86344 68869 86379 68897
rect 86407 68869 86441 68897
rect 86469 68869 86504 68897
rect 86344 68835 86504 68869
rect 86344 68807 86379 68835
rect 86407 68807 86441 68835
rect 86469 68807 86504 68835
rect 86344 68773 86504 68807
rect 86344 68745 86379 68773
rect 86407 68745 86441 68773
rect 86469 68745 86504 68773
rect 86344 68728 86504 68745
rect 101704 68959 101864 68976
rect 101704 68931 101739 68959
rect 101767 68931 101801 68959
rect 101829 68931 101864 68959
rect 101704 68897 101864 68931
rect 101704 68869 101739 68897
rect 101767 68869 101801 68897
rect 101829 68869 101864 68897
rect 101704 68835 101864 68869
rect 101704 68807 101739 68835
rect 101767 68807 101801 68835
rect 101829 68807 101864 68835
rect 101704 68773 101864 68807
rect 101704 68745 101739 68773
rect 101767 68745 101801 68773
rect 101829 68745 101864 68773
rect 101704 68728 101864 68745
rect 117064 68959 117224 68976
rect 117064 68931 117099 68959
rect 117127 68931 117161 68959
rect 117189 68931 117224 68959
rect 117064 68897 117224 68931
rect 117064 68869 117099 68897
rect 117127 68869 117161 68897
rect 117189 68869 117224 68897
rect 117064 68835 117224 68869
rect 117064 68807 117099 68835
rect 117127 68807 117161 68835
rect 117189 68807 117224 68835
rect 117064 68773 117224 68807
rect 117064 68745 117099 68773
rect 117127 68745 117161 68773
rect 117189 68745 117224 68773
rect 117064 68728 117224 68745
rect 132424 68959 132584 68976
rect 132424 68931 132459 68959
rect 132487 68931 132521 68959
rect 132549 68931 132584 68959
rect 132424 68897 132584 68931
rect 132424 68869 132459 68897
rect 132487 68869 132521 68897
rect 132549 68869 132584 68897
rect 132424 68835 132584 68869
rect 132424 68807 132459 68835
rect 132487 68807 132521 68835
rect 132549 68807 132584 68835
rect 132424 68773 132584 68807
rect 132424 68745 132459 68773
rect 132487 68745 132521 68773
rect 132549 68745 132584 68773
rect 132424 68728 132584 68745
rect 147784 68959 147944 68976
rect 147784 68931 147819 68959
rect 147847 68931 147881 68959
rect 147909 68931 147944 68959
rect 147784 68897 147944 68931
rect 147784 68869 147819 68897
rect 147847 68869 147881 68897
rect 147909 68869 147944 68897
rect 147784 68835 147944 68869
rect 147784 68807 147819 68835
rect 147847 68807 147881 68835
rect 147909 68807 147944 68835
rect 147784 68773 147944 68807
rect 147784 68745 147819 68773
rect 147847 68745 147881 68773
rect 147909 68745 147944 68773
rect 147784 68728 147944 68745
rect 163144 68959 163304 68976
rect 163144 68931 163179 68959
rect 163207 68931 163241 68959
rect 163269 68931 163304 68959
rect 163144 68897 163304 68931
rect 163144 68869 163179 68897
rect 163207 68869 163241 68897
rect 163269 68869 163304 68897
rect 163144 68835 163304 68869
rect 163144 68807 163179 68835
rect 163207 68807 163241 68835
rect 163269 68807 163304 68835
rect 163144 68773 163304 68807
rect 163144 68745 163179 68773
rect 163207 68745 163241 68773
rect 163269 68745 163304 68773
rect 163144 68728 163304 68745
rect 178504 68959 178664 68976
rect 178504 68931 178539 68959
rect 178567 68931 178601 68959
rect 178629 68931 178664 68959
rect 178504 68897 178664 68931
rect 178504 68869 178539 68897
rect 178567 68869 178601 68897
rect 178629 68869 178664 68897
rect 178504 68835 178664 68869
rect 178504 68807 178539 68835
rect 178567 68807 178601 68835
rect 178629 68807 178664 68835
rect 178504 68773 178664 68807
rect 178504 68745 178539 68773
rect 178567 68745 178601 68773
rect 178629 68745 178664 68773
rect 178504 68728 178664 68745
rect 193864 68959 194024 68976
rect 193864 68931 193899 68959
rect 193927 68931 193961 68959
rect 193989 68931 194024 68959
rect 193864 68897 194024 68931
rect 193864 68869 193899 68897
rect 193927 68869 193961 68897
rect 193989 68869 194024 68897
rect 193864 68835 194024 68869
rect 193864 68807 193899 68835
rect 193927 68807 193961 68835
rect 193989 68807 194024 68835
rect 193864 68773 194024 68807
rect 193864 68745 193899 68773
rect 193927 68745 193961 68773
rect 193989 68745 194024 68773
rect 193864 68728 194024 68745
rect 209224 68959 209384 68976
rect 209224 68931 209259 68959
rect 209287 68931 209321 68959
rect 209349 68931 209384 68959
rect 209224 68897 209384 68931
rect 209224 68869 209259 68897
rect 209287 68869 209321 68897
rect 209349 68869 209384 68897
rect 209224 68835 209384 68869
rect 209224 68807 209259 68835
rect 209287 68807 209321 68835
rect 209349 68807 209384 68835
rect 209224 68773 209384 68807
rect 209224 68745 209259 68773
rect 209287 68745 209321 68773
rect 209349 68745 209384 68773
rect 209224 68728 209384 68745
rect 224584 68959 224744 68976
rect 224584 68931 224619 68959
rect 224647 68931 224681 68959
rect 224709 68931 224744 68959
rect 224584 68897 224744 68931
rect 224584 68869 224619 68897
rect 224647 68869 224681 68897
rect 224709 68869 224744 68897
rect 224584 68835 224744 68869
rect 224584 68807 224619 68835
rect 224647 68807 224681 68835
rect 224709 68807 224744 68835
rect 224584 68773 224744 68807
rect 224584 68745 224619 68773
rect 224647 68745 224681 68773
rect 224709 68745 224744 68773
rect 224584 68728 224744 68745
rect 239944 68959 240104 68976
rect 239944 68931 239979 68959
rect 240007 68931 240041 68959
rect 240069 68931 240104 68959
rect 239944 68897 240104 68931
rect 239944 68869 239979 68897
rect 240007 68869 240041 68897
rect 240069 68869 240104 68897
rect 239944 68835 240104 68869
rect 239944 68807 239979 68835
rect 240007 68807 240041 68835
rect 240069 68807 240104 68835
rect 239944 68773 240104 68807
rect 239944 68745 239979 68773
rect 240007 68745 240041 68773
rect 240069 68745 240104 68773
rect 239944 68728 240104 68745
rect 32584 65959 32744 65976
rect 32584 65931 32619 65959
rect 32647 65931 32681 65959
rect 32709 65931 32744 65959
rect 32584 65897 32744 65931
rect 32584 65869 32619 65897
rect 32647 65869 32681 65897
rect 32709 65869 32744 65897
rect 32584 65835 32744 65869
rect 32584 65807 32619 65835
rect 32647 65807 32681 65835
rect 32709 65807 32744 65835
rect 32584 65773 32744 65807
rect 32584 65745 32619 65773
rect 32647 65745 32681 65773
rect 32709 65745 32744 65773
rect 32584 65728 32744 65745
rect 47944 65959 48104 65976
rect 47944 65931 47979 65959
rect 48007 65931 48041 65959
rect 48069 65931 48104 65959
rect 47944 65897 48104 65931
rect 47944 65869 47979 65897
rect 48007 65869 48041 65897
rect 48069 65869 48104 65897
rect 47944 65835 48104 65869
rect 47944 65807 47979 65835
rect 48007 65807 48041 65835
rect 48069 65807 48104 65835
rect 47944 65773 48104 65807
rect 47944 65745 47979 65773
rect 48007 65745 48041 65773
rect 48069 65745 48104 65773
rect 47944 65728 48104 65745
rect 63304 65959 63464 65976
rect 63304 65931 63339 65959
rect 63367 65931 63401 65959
rect 63429 65931 63464 65959
rect 63304 65897 63464 65931
rect 63304 65869 63339 65897
rect 63367 65869 63401 65897
rect 63429 65869 63464 65897
rect 63304 65835 63464 65869
rect 63304 65807 63339 65835
rect 63367 65807 63401 65835
rect 63429 65807 63464 65835
rect 63304 65773 63464 65807
rect 63304 65745 63339 65773
rect 63367 65745 63401 65773
rect 63429 65745 63464 65773
rect 63304 65728 63464 65745
rect 78664 65959 78824 65976
rect 78664 65931 78699 65959
rect 78727 65931 78761 65959
rect 78789 65931 78824 65959
rect 78664 65897 78824 65931
rect 78664 65869 78699 65897
rect 78727 65869 78761 65897
rect 78789 65869 78824 65897
rect 78664 65835 78824 65869
rect 78664 65807 78699 65835
rect 78727 65807 78761 65835
rect 78789 65807 78824 65835
rect 78664 65773 78824 65807
rect 78664 65745 78699 65773
rect 78727 65745 78761 65773
rect 78789 65745 78824 65773
rect 78664 65728 78824 65745
rect 94024 65959 94184 65976
rect 94024 65931 94059 65959
rect 94087 65931 94121 65959
rect 94149 65931 94184 65959
rect 94024 65897 94184 65931
rect 94024 65869 94059 65897
rect 94087 65869 94121 65897
rect 94149 65869 94184 65897
rect 94024 65835 94184 65869
rect 94024 65807 94059 65835
rect 94087 65807 94121 65835
rect 94149 65807 94184 65835
rect 94024 65773 94184 65807
rect 94024 65745 94059 65773
rect 94087 65745 94121 65773
rect 94149 65745 94184 65773
rect 94024 65728 94184 65745
rect 109384 65959 109544 65976
rect 109384 65931 109419 65959
rect 109447 65931 109481 65959
rect 109509 65931 109544 65959
rect 109384 65897 109544 65931
rect 109384 65869 109419 65897
rect 109447 65869 109481 65897
rect 109509 65869 109544 65897
rect 109384 65835 109544 65869
rect 109384 65807 109419 65835
rect 109447 65807 109481 65835
rect 109509 65807 109544 65835
rect 109384 65773 109544 65807
rect 109384 65745 109419 65773
rect 109447 65745 109481 65773
rect 109509 65745 109544 65773
rect 109384 65728 109544 65745
rect 124744 65959 124904 65976
rect 124744 65931 124779 65959
rect 124807 65931 124841 65959
rect 124869 65931 124904 65959
rect 124744 65897 124904 65931
rect 124744 65869 124779 65897
rect 124807 65869 124841 65897
rect 124869 65869 124904 65897
rect 124744 65835 124904 65869
rect 124744 65807 124779 65835
rect 124807 65807 124841 65835
rect 124869 65807 124904 65835
rect 124744 65773 124904 65807
rect 124744 65745 124779 65773
rect 124807 65745 124841 65773
rect 124869 65745 124904 65773
rect 124744 65728 124904 65745
rect 140104 65959 140264 65976
rect 140104 65931 140139 65959
rect 140167 65931 140201 65959
rect 140229 65931 140264 65959
rect 140104 65897 140264 65931
rect 140104 65869 140139 65897
rect 140167 65869 140201 65897
rect 140229 65869 140264 65897
rect 140104 65835 140264 65869
rect 140104 65807 140139 65835
rect 140167 65807 140201 65835
rect 140229 65807 140264 65835
rect 140104 65773 140264 65807
rect 140104 65745 140139 65773
rect 140167 65745 140201 65773
rect 140229 65745 140264 65773
rect 140104 65728 140264 65745
rect 155464 65959 155624 65976
rect 155464 65931 155499 65959
rect 155527 65931 155561 65959
rect 155589 65931 155624 65959
rect 155464 65897 155624 65931
rect 155464 65869 155499 65897
rect 155527 65869 155561 65897
rect 155589 65869 155624 65897
rect 155464 65835 155624 65869
rect 155464 65807 155499 65835
rect 155527 65807 155561 65835
rect 155589 65807 155624 65835
rect 155464 65773 155624 65807
rect 155464 65745 155499 65773
rect 155527 65745 155561 65773
rect 155589 65745 155624 65773
rect 155464 65728 155624 65745
rect 170824 65959 170984 65976
rect 170824 65931 170859 65959
rect 170887 65931 170921 65959
rect 170949 65931 170984 65959
rect 170824 65897 170984 65931
rect 170824 65869 170859 65897
rect 170887 65869 170921 65897
rect 170949 65869 170984 65897
rect 170824 65835 170984 65869
rect 170824 65807 170859 65835
rect 170887 65807 170921 65835
rect 170949 65807 170984 65835
rect 170824 65773 170984 65807
rect 170824 65745 170859 65773
rect 170887 65745 170921 65773
rect 170949 65745 170984 65773
rect 170824 65728 170984 65745
rect 186184 65959 186344 65976
rect 186184 65931 186219 65959
rect 186247 65931 186281 65959
rect 186309 65931 186344 65959
rect 186184 65897 186344 65931
rect 186184 65869 186219 65897
rect 186247 65869 186281 65897
rect 186309 65869 186344 65897
rect 186184 65835 186344 65869
rect 186184 65807 186219 65835
rect 186247 65807 186281 65835
rect 186309 65807 186344 65835
rect 186184 65773 186344 65807
rect 186184 65745 186219 65773
rect 186247 65745 186281 65773
rect 186309 65745 186344 65773
rect 186184 65728 186344 65745
rect 201544 65959 201704 65976
rect 201544 65931 201579 65959
rect 201607 65931 201641 65959
rect 201669 65931 201704 65959
rect 201544 65897 201704 65931
rect 201544 65869 201579 65897
rect 201607 65869 201641 65897
rect 201669 65869 201704 65897
rect 201544 65835 201704 65869
rect 201544 65807 201579 65835
rect 201607 65807 201641 65835
rect 201669 65807 201704 65835
rect 201544 65773 201704 65807
rect 201544 65745 201579 65773
rect 201607 65745 201641 65773
rect 201669 65745 201704 65773
rect 201544 65728 201704 65745
rect 216904 65959 217064 65976
rect 216904 65931 216939 65959
rect 216967 65931 217001 65959
rect 217029 65931 217064 65959
rect 216904 65897 217064 65931
rect 216904 65869 216939 65897
rect 216967 65869 217001 65897
rect 217029 65869 217064 65897
rect 216904 65835 217064 65869
rect 216904 65807 216939 65835
rect 216967 65807 217001 65835
rect 217029 65807 217064 65835
rect 216904 65773 217064 65807
rect 216904 65745 216939 65773
rect 216967 65745 217001 65773
rect 217029 65745 217064 65773
rect 216904 65728 217064 65745
rect 232264 65959 232424 65976
rect 232264 65931 232299 65959
rect 232327 65931 232361 65959
rect 232389 65931 232424 65959
rect 232264 65897 232424 65931
rect 232264 65869 232299 65897
rect 232327 65869 232361 65897
rect 232389 65869 232424 65897
rect 232264 65835 232424 65869
rect 232264 65807 232299 65835
rect 232327 65807 232361 65835
rect 232389 65807 232424 65835
rect 232264 65773 232424 65807
rect 232264 65745 232299 65773
rect 232327 65745 232361 65773
rect 232389 65745 232424 65773
rect 232264 65728 232424 65745
rect 247624 65959 247784 65976
rect 247624 65931 247659 65959
rect 247687 65931 247721 65959
rect 247749 65931 247784 65959
rect 247624 65897 247784 65931
rect 247624 65869 247659 65897
rect 247687 65869 247721 65897
rect 247749 65869 247784 65897
rect 247624 65835 247784 65869
rect 247624 65807 247659 65835
rect 247687 65807 247721 65835
rect 247749 65807 247784 65835
rect 247624 65773 247784 65807
rect 247624 65745 247659 65773
rect 247687 65745 247721 65773
rect 247749 65745 247784 65773
rect 247624 65728 247784 65745
rect 254529 65959 254839 74745
rect 254529 65931 254577 65959
rect 254605 65931 254639 65959
rect 254667 65931 254701 65959
rect 254729 65931 254763 65959
rect 254791 65931 254839 65959
rect 254529 65897 254839 65931
rect 254529 65869 254577 65897
rect 254605 65869 254639 65897
rect 254667 65869 254701 65897
rect 254729 65869 254763 65897
rect 254791 65869 254839 65897
rect 254529 65835 254839 65869
rect 254529 65807 254577 65835
rect 254605 65807 254639 65835
rect 254667 65807 254701 65835
rect 254729 65807 254763 65835
rect 254791 65807 254839 65835
rect 254529 65773 254839 65807
rect 254529 65745 254577 65773
rect 254605 65745 254639 65773
rect 254667 65745 254701 65773
rect 254729 65745 254763 65773
rect 254791 65745 254839 65773
rect 31389 59931 31437 59959
rect 31465 59931 31499 59959
rect 31527 59931 31561 59959
rect 31589 59931 31623 59959
rect 31651 59931 31699 59959
rect 31389 59897 31699 59931
rect 31389 59869 31437 59897
rect 31465 59869 31499 59897
rect 31527 59869 31561 59897
rect 31589 59869 31623 59897
rect 31651 59869 31699 59897
rect 31389 59835 31699 59869
rect 31389 59807 31437 59835
rect 31465 59807 31499 59835
rect 31527 59807 31561 59835
rect 31589 59807 31623 59835
rect 31651 59807 31699 59835
rect 31389 59773 31699 59807
rect 31389 59745 31437 59773
rect 31465 59745 31499 59773
rect 31527 59745 31561 59773
rect 31589 59745 31623 59773
rect 31651 59745 31699 59773
rect 31389 50959 31699 59745
rect 40264 59959 40424 59976
rect 40264 59931 40299 59959
rect 40327 59931 40361 59959
rect 40389 59931 40424 59959
rect 40264 59897 40424 59931
rect 40264 59869 40299 59897
rect 40327 59869 40361 59897
rect 40389 59869 40424 59897
rect 40264 59835 40424 59869
rect 40264 59807 40299 59835
rect 40327 59807 40361 59835
rect 40389 59807 40424 59835
rect 40264 59773 40424 59807
rect 40264 59745 40299 59773
rect 40327 59745 40361 59773
rect 40389 59745 40424 59773
rect 40264 59728 40424 59745
rect 55624 59959 55784 59976
rect 55624 59931 55659 59959
rect 55687 59931 55721 59959
rect 55749 59931 55784 59959
rect 55624 59897 55784 59931
rect 55624 59869 55659 59897
rect 55687 59869 55721 59897
rect 55749 59869 55784 59897
rect 55624 59835 55784 59869
rect 55624 59807 55659 59835
rect 55687 59807 55721 59835
rect 55749 59807 55784 59835
rect 55624 59773 55784 59807
rect 55624 59745 55659 59773
rect 55687 59745 55721 59773
rect 55749 59745 55784 59773
rect 55624 59728 55784 59745
rect 70984 59959 71144 59976
rect 70984 59931 71019 59959
rect 71047 59931 71081 59959
rect 71109 59931 71144 59959
rect 70984 59897 71144 59931
rect 70984 59869 71019 59897
rect 71047 59869 71081 59897
rect 71109 59869 71144 59897
rect 70984 59835 71144 59869
rect 70984 59807 71019 59835
rect 71047 59807 71081 59835
rect 71109 59807 71144 59835
rect 70984 59773 71144 59807
rect 70984 59745 71019 59773
rect 71047 59745 71081 59773
rect 71109 59745 71144 59773
rect 70984 59728 71144 59745
rect 86344 59959 86504 59976
rect 86344 59931 86379 59959
rect 86407 59931 86441 59959
rect 86469 59931 86504 59959
rect 86344 59897 86504 59931
rect 86344 59869 86379 59897
rect 86407 59869 86441 59897
rect 86469 59869 86504 59897
rect 86344 59835 86504 59869
rect 86344 59807 86379 59835
rect 86407 59807 86441 59835
rect 86469 59807 86504 59835
rect 86344 59773 86504 59807
rect 86344 59745 86379 59773
rect 86407 59745 86441 59773
rect 86469 59745 86504 59773
rect 86344 59728 86504 59745
rect 101704 59959 101864 59976
rect 101704 59931 101739 59959
rect 101767 59931 101801 59959
rect 101829 59931 101864 59959
rect 101704 59897 101864 59931
rect 101704 59869 101739 59897
rect 101767 59869 101801 59897
rect 101829 59869 101864 59897
rect 101704 59835 101864 59869
rect 101704 59807 101739 59835
rect 101767 59807 101801 59835
rect 101829 59807 101864 59835
rect 101704 59773 101864 59807
rect 101704 59745 101739 59773
rect 101767 59745 101801 59773
rect 101829 59745 101864 59773
rect 101704 59728 101864 59745
rect 117064 59959 117224 59976
rect 117064 59931 117099 59959
rect 117127 59931 117161 59959
rect 117189 59931 117224 59959
rect 117064 59897 117224 59931
rect 117064 59869 117099 59897
rect 117127 59869 117161 59897
rect 117189 59869 117224 59897
rect 117064 59835 117224 59869
rect 117064 59807 117099 59835
rect 117127 59807 117161 59835
rect 117189 59807 117224 59835
rect 117064 59773 117224 59807
rect 117064 59745 117099 59773
rect 117127 59745 117161 59773
rect 117189 59745 117224 59773
rect 117064 59728 117224 59745
rect 132424 59959 132584 59976
rect 132424 59931 132459 59959
rect 132487 59931 132521 59959
rect 132549 59931 132584 59959
rect 132424 59897 132584 59931
rect 132424 59869 132459 59897
rect 132487 59869 132521 59897
rect 132549 59869 132584 59897
rect 132424 59835 132584 59869
rect 132424 59807 132459 59835
rect 132487 59807 132521 59835
rect 132549 59807 132584 59835
rect 132424 59773 132584 59807
rect 132424 59745 132459 59773
rect 132487 59745 132521 59773
rect 132549 59745 132584 59773
rect 132424 59728 132584 59745
rect 147784 59959 147944 59976
rect 147784 59931 147819 59959
rect 147847 59931 147881 59959
rect 147909 59931 147944 59959
rect 147784 59897 147944 59931
rect 147784 59869 147819 59897
rect 147847 59869 147881 59897
rect 147909 59869 147944 59897
rect 147784 59835 147944 59869
rect 147784 59807 147819 59835
rect 147847 59807 147881 59835
rect 147909 59807 147944 59835
rect 147784 59773 147944 59807
rect 147784 59745 147819 59773
rect 147847 59745 147881 59773
rect 147909 59745 147944 59773
rect 147784 59728 147944 59745
rect 163144 59959 163304 59976
rect 163144 59931 163179 59959
rect 163207 59931 163241 59959
rect 163269 59931 163304 59959
rect 163144 59897 163304 59931
rect 163144 59869 163179 59897
rect 163207 59869 163241 59897
rect 163269 59869 163304 59897
rect 163144 59835 163304 59869
rect 163144 59807 163179 59835
rect 163207 59807 163241 59835
rect 163269 59807 163304 59835
rect 163144 59773 163304 59807
rect 163144 59745 163179 59773
rect 163207 59745 163241 59773
rect 163269 59745 163304 59773
rect 163144 59728 163304 59745
rect 178504 59959 178664 59976
rect 178504 59931 178539 59959
rect 178567 59931 178601 59959
rect 178629 59931 178664 59959
rect 178504 59897 178664 59931
rect 178504 59869 178539 59897
rect 178567 59869 178601 59897
rect 178629 59869 178664 59897
rect 178504 59835 178664 59869
rect 178504 59807 178539 59835
rect 178567 59807 178601 59835
rect 178629 59807 178664 59835
rect 178504 59773 178664 59807
rect 178504 59745 178539 59773
rect 178567 59745 178601 59773
rect 178629 59745 178664 59773
rect 178504 59728 178664 59745
rect 193864 59959 194024 59976
rect 193864 59931 193899 59959
rect 193927 59931 193961 59959
rect 193989 59931 194024 59959
rect 193864 59897 194024 59931
rect 193864 59869 193899 59897
rect 193927 59869 193961 59897
rect 193989 59869 194024 59897
rect 193864 59835 194024 59869
rect 193864 59807 193899 59835
rect 193927 59807 193961 59835
rect 193989 59807 194024 59835
rect 193864 59773 194024 59807
rect 193864 59745 193899 59773
rect 193927 59745 193961 59773
rect 193989 59745 194024 59773
rect 193864 59728 194024 59745
rect 209224 59959 209384 59976
rect 209224 59931 209259 59959
rect 209287 59931 209321 59959
rect 209349 59931 209384 59959
rect 209224 59897 209384 59931
rect 209224 59869 209259 59897
rect 209287 59869 209321 59897
rect 209349 59869 209384 59897
rect 209224 59835 209384 59869
rect 209224 59807 209259 59835
rect 209287 59807 209321 59835
rect 209349 59807 209384 59835
rect 209224 59773 209384 59807
rect 209224 59745 209259 59773
rect 209287 59745 209321 59773
rect 209349 59745 209384 59773
rect 209224 59728 209384 59745
rect 224584 59959 224744 59976
rect 224584 59931 224619 59959
rect 224647 59931 224681 59959
rect 224709 59931 224744 59959
rect 224584 59897 224744 59931
rect 224584 59869 224619 59897
rect 224647 59869 224681 59897
rect 224709 59869 224744 59897
rect 224584 59835 224744 59869
rect 224584 59807 224619 59835
rect 224647 59807 224681 59835
rect 224709 59807 224744 59835
rect 224584 59773 224744 59807
rect 224584 59745 224619 59773
rect 224647 59745 224681 59773
rect 224709 59745 224744 59773
rect 224584 59728 224744 59745
rect 239944 59959 240104 59976
rect 239944 59931 239979 59959
rect 240007 59931 240041 59959
rect 240069 59931 240104 59959
rect 239944 59897 240104 59931
rect 239944 59869 239979 59897
rect 240007 59869 240041 59897
rect 240069 59869 240104 59897
rect 239944 59835 240104 59869
rect 239944 59807 239979 59835
rect 240007 59807 240041 59835
rect 240069 59807 240104 59835
rect 239944 59773 240104 59807
rect 239944 59745 239979 59773
rect 240007 59745 240041 59773
rect 240069 59745 240104 59773
rect 239944 59728 240104 59745
rect 32584 56959 32744 56976
rect 32584 56931 32619 56959
rect 32647 56931 32681 56959
rect 32709 56931 32744 56959
rect 32584 56897 32744 56931
rect 32584 56869 32619 56897
rect 32647 56869 32681 56897
rect 32709 56869 32744 56897
rect 32584 56835 32744 56869
rect 32584 56807 32619 56835
rect 32647 56807 32681 56835
rect 32709 56807 32744 56835
rect 32584 56773 32744 56807
rect 32584 56745 32619 56773
rect 32647 56745 32681 56773
rect 32709 56745 32744 56773
rect 32584 56728 32744 56745
rect 47944 56959 48104 56976
rect 47944 56931 47979 56959
rect 48007 56931 48041 56959
rect 48069 56931 48104 56959
rect 47944 56897 48104 56931
rect 47944 56869 47979 56897
rect 48007 56869 48041 56897
rect 48069 56869 48104 56897
rect 47944 56835 48104 56869
rect 47944 56807 47979 56835
rect 48007 56807 48041 56835
rect 48069 56807 48104 56835
rect 47944 56773 48104 56807
rect 47944 56745 47979 56773
rect 48007 56745 48041 56773
rect 48069 56745 48104 56773
rect 47944 56728 48104 56745
rect 63304 56959 63464 56976
rect 63304 56931 63339 56959
rect 63367 56931 63401 56959
rect 63429 56931 63464 56959
rect 63304 56897 63464 56931
rect 63304 56869 63339 56897
rect 63367 56869 63401 56897
rect 63429 56869 63464 56897
rect 63304 56835 63464 56869
rect 63304 56807 63339 56835
rect 63367 56807 63401 56835
rect 63429 56807 63464 56835
rect 63304 56773 63464 56807
rect 63304 56745 63339 56773
rect 63367 56745 63401 56773
rect 63429 56745 63464 56773
rect 63304 56728 63464 56745
rect 78664 56959 78824 56976
rect 78664 56931 78699 56959
rect 78727 56931 78761 56959
rect 78789 56931 78824 56959
rect 78664 56897 78824 56931
rect 78664 56869 78699 56897
rect 78727 56869 78761 56897
rect 78789 56869 78824 56897
rect 78664 56835 78824 56869
rect 78664 56807 78699 56835
rect 78727 56807 78761 56835
rect 78789 56807 78824 56835
rect 78664 56773 78824 56807
rect 78664 56745 78699 56773
rect 78727 56745 78761 56773
rect 78789 56745 78824 56773
rect 78664 56728 78824 56745
rect 94024 56959 94184 56976
rect 94024 56931 94059 56959
rect 94087 56931 94121 56959
rect 94149 56931 94184 56959
rect 94024 56897 94184 56931
rect 94024 56869 94059 56897
rect 94087 56869 94121 56897
rect 94149 56869 94184 56897
rect 94024 56835 94184 56869
rect 94024 56807 94059 56835
rect 94087 56807 94121 56835
rect 94149 56807 94184 56835
rect 94024 56773 94184 56807
rect 94024 56745 94059 56773
rect 94087 56745 94121 56773
rect 94149 56745 94184 56773
rect 94024 56728 94184 56745
rect 109384 56959 109544 56976
rect 109384 56931 109419 56959
rect 109447 56931 109481 56959
rect 109509 56931 109544 56959
rect 109384 56897 109544 56931
rect 109384 56869 109419 56897
rect 109447 56869 109481 56897
rect 109509 56869 109544 56897
rect 109384 56835 109544 56869
rect 109384 56807 109419 56835
rect 109447 56807 109481 56835
rect 109509 56807 109544 56835
rect 109384 56773 109544 56807
rect 109384 56745 109419 56773
rect 109447 56745 109481 56773
rect 109509 56745 109544 56773
rect 109384 56728 109544 56745
rect 124744 56959 124904 56976
rect 124744 56931 124779 56959
rect 124807 56931 124841 56959
rect 124869 56931 124904 56959
rect 124744 56897 124904 56931
rect 124744 56869 124779 56897
rect 124807 56869 124841 56897
rect 124869 56869 124904 56897
rect 124744 56835 124904 56869
rect 124744 56807 124779 56835
rect 124807 56807 124841 56835
rect 124869 56807 124904 56835
rect 124744 56773 124904 56807
rect 124744 56745 124779 56773
rect 124807 56745 124841 56773
rect 124869 56745 124904 56773
rect 124744 56728 124904 56745
rect 140104 56959 140264 56976
rect 140104 56931 140139 56959
rect 140167 56931 140201 56959
rect 140229 56931 140264 56959
rect 140104 56897 140264 56931
rect 140104 56869 140139 56897
rect 140167 56869 140201 56897
rect 140229 56869 140264 56897
rect 140104 56835 140264 56869
rect 140104 56807 140139 56835
rect 140167 56807 140201 56835
rect 140229 56807 140264 56835
rect 140104 56773 140264 56807
rect 140104 56745 140139 56773
rect 140167 56745 140201 56773
rect 140229 56745 140264 56773
rect 140104 56728 140264 56745
rect 155464 56959 155624 56976
rect 155464 56931 155499 56959
rect 155527 56931 155561 56959
rect 155589 56931 155624 56959
rect 155464 56897 155624 56931
rect 155464 56869 155499 56897
rect 155527 56869 155561 56897
rect 155589 56869 155624 56897
rect 155464 56835 155624 56869
rect 155464 56807 155499 56835
rect 155527 56807 155561 56835
rect 155589 56807 155624 56835
rect 155464 56773 155624 56807
rect 155464 56745 155499 56773
rect 155527 56745 155561 56773
rect 155589 56745 155624 56773
rect 155464 56728 155624 56745
rect 170824 56959 170984 56976
rect 170824 56931 170859 56959
rect 170887 56931 170921 56959
rect 170949 56931 170984 56959
rect 170824 56897 170984 56931
rect 170824 56869 170859 56897
rect 170887 56869 170921 56897
rect 170949 56869 170984 56897
rect 170824 56835 170984 56869
rect 170824 56807 170859 56835
rect 170887 56807 170921 56835
rect 170949 56807 170984 56835
rect 170824 56773 170984 56807
rect 170824 56745 170859 56773
rect 170887 56745 170921 56773
rect 170949 56745 170984 56773
rect 170824 56728 170984 56745
rect 186184 56959 186344 56976
rect 186184 56931 186219 56959
rect 186247 56931 186281 56959
rect 186309 56931 186344 56959
rect 186184 56897 186344 56931
rect 186184 56869 186219 56897
rect 186247 56869 186281 56897
rect 186309 56869 186344 56897
rect 186184 56835 186344 56869
rect 186184 56807 186219 56835
rect 186247 56807 186281 56835
rect 186309 56807 186344 56835
rect 186184 56773 186344 56807
rect 186184 56745 186219 56773
rect 186247 56745 186281 56773
rect 186309 56745 186344 56773
rect 186184 56728 186344 56745
rect 201544 56959 201704 56976
rect 201544 56931 201579 56959
rect 201607 56931 201641 56959
rect 201669 56931 201704 56959
rect 201544 56897 201704 56931
rect 201544 56869 201579 56897
rect 201607 56869 201641 56897
rect 201669 56869 201704 56897
rect 201544 56835 201704 56869
rect 201544 56807 201579 56835
rect 201607 56807 201641 56835
rect 201669 56807 201704 56835
rect 201544 56773 201704 56807
rect 201544 56745 201579 56773
rect 201607 56745 201641 56773
rect 201669 56745 201704 56773
rect 201544 56728 201704 56745
rect 216904 56959 217064 56976
rect 216904 56931 216939 56959
rect 216967 56931 217001 56959
rect 217029 56931 217064 56959
rect 216904 56897 217064 56931
rect 216904 56869 216939 56897
rect 216967 56869 217001 56897
rect 217029 56869 217064 56897
rect 216904 56835 217064 56869
rect 216904 56807 216939 56835
rect 216967 56807 217001 56835
rect 217029 56807 217064 56835
rect 216904 56773 217064 56807
rect 216904 56745 216939 56773
rect 216967 56745 217001 56773
rect 217029 56745 217064 56773
rect 216904 56728 217064 56745
rect 232264 56959 232424 56976
rect 232264 56931 232299 56959
rect 232327 56931 232361 56959
rect 232389 56931 232424 56959
rect 232264 56897 232424 56931
rect 232264 56869 232299 56897
rect 232327 56869 232361 56897
rect 232389 56869 232424 56897
rect 232264 56835 232424 56869
rect 232264 56807 232299 56835
rect 232327 56807 232361 56835
rect 232389 56807 232424 56835
rect 232264 56773 232424 56807
rect 232264 56745 232299 56773
rect 232327 56745 232361 56773
rect 232389 56745 232424 56773
rect 232264 56728 232424 56745
rect 247624 56959 247784 56976
rect 247624 56931 247659 56959
rect 247687 56931 247721 56959
rect 247749 56931 247784 56959
rect 247624 56897 247784 56931
rect 247624 56869 247659 56897
rect 247687 56869 247721 56897
rect 247749 56869 247784 56897
rect 247624 56835 247784 56869
rect 247624 56807 247659 56835
rect 247687 56807 247721 56835
rect 247749 56807 247784 56835
rect 247624 56773 247784 56807
rect 247624 56745 247659 56773
rect 247687 56745 247721 56773
rect 247749 56745 247784 56773
rect 247624 56728 247784 56745
rect 254529 56959 254839 65745
rect 254529 56931 254577 56959
rect 254605 56931 254639 56959
rect 254667 56931 254701 56959
rect 254729 56931 254763 56959
rect 254791 56931 254839 56959
rect 254529 56897 254839 56931
rect 254529 56869 254577 56897
rect 254605 56869 254639 56897
rect 254667 56869 254701 56897
rect 254729 56869 254763 56897
rect 254791 56869 254839 56897
rect 254529 56835 254839 56869
rect 254529 56807 254577 56835
rect 254605 56807 254639 56835
rect 254667 56807 254701 56835
rect 254729 56807 254763 56835
rect 254791 56807 254839 56835
rect 254529 56773 254839 56807
rect 254529 56745 254577 56773
rect 254605 56745 254639 56773
rect 254667 56745 254701 56773
rect 254729 56745 254763 56773
rect 254791 56745 254839 56773
rect 31389 50931 31437 50959
rect 31465 50931 31499 50959
rect 31527 50931 31561 50959
rect 31589 50931 31623 50959
rect 31651 50931 31699 50959
rect 31389 50897 31699 50931
rect 31389 50869 31437 50897
rect 31465 50869 31499 50897
rect 31527 50869 31561 50897
rect 31589 50869 31623 50897
rect 31651 50869 31699 50897
rect 31389 50835 31699 50869
rect 31389 50807 31437 50835
rect 31465 50807 31499 50835
rect 31527 50807 31561 50835
rect 31589 50807 31623 50835
rect 31651 50807 31699 50835
rect 31389 50773 31699 50807
rect 31389 50745 31437 50773
rect 31465 50745 31499 50773
rect 31527 50745 31561 50773
rect 31589 50745 31623 50773
rect 31651 50745 31699 50773
rect 31389 41959 31699 50745
rect 40264 50959 40424 50976
rect 40264 50931 40299 50959
rect 40327 50931 40361 50959
rect 40389 50931 40424 50959
rect 40264 50897 40424 50931
rect 40264 50869 40299 50897
rect 40327 50869 40361 50897
rect 40389 50869 40424 50897
rect 40264 50835 40424 50869
rect 40264 50807 40299 50835
rect 40327 50807 40361 50835
rect 40389 50807 40424 50835
rect 40264 50773 40424 50807
rect 40264 50745 40299 50773
rect 40327 50745 40361 50773
rect 40389 50745 40424 50773
rect 40264 50728 40424 50745
rect 55624 50959 55784 50976
rect 55624 50931 55659 50959
rect 55687 50931 55721 50959
rect 55749 50931 55784 50959
rect 55624 50897 55784 50931
rect 55624 50869 55659 50897
rect 55687 50869 55721 50897
rect 55749 50869 55784 50897
rect 55624 50835 55784 50869
rect 55624 50807 55659 50835
rect 55687 50807 55721 50835
rect 55749 50807 55784 50835
rect 55624 50773 55784 50807
rect 55624 50745 55659 50773
rect 55687 50745 55721 50773
rect 55749 50745 55784 50773
rect 55624 50728 55784 50745
rect 70984 50959 71144 50976
rect 70984 50931 71019 50959
rect 71047 50931 71081 50959
rect 71109 50931 71144 50959
rect 70984 50897 71144 50931
rect 70984 50869 71019 50897
rect 71047 50869 71081 50897
rect 71109 50869 71144 50897
rect 70984 50835 71144 50869
rect 70984 50807 71019 50835
rect 71047 50807 71081 50835
rect 71109 50807 71144 50835
rect 70984 50773 71144 50807
rect 70984 50745 71019 50773
rect 71047 50745 71081 50773
rect 71109 50745 71144 50773
rect 70984 50728 71144 50745
rect 86344 50959 86504 50976
rect 86344 50931 86379 50959
rect 86407 50931 86441 50959
rect 86469 50931 86504 50959
rect 86344 50897 86504 50931
rect 86344 50869 86379 50897
rect 86407 50869 86441 50897
rect 86469 50869 86504 50897
rect 86344 50835 86504 50869
rect 86344 50807 86379 50835
rect 86407 50807 86441 50835
rect 86469 50807 86504 50835
rect 86344 50773 86504 50807
rect 86344 50745 86379 50773
rect 86407 50745 86441 50773
rect 86469 50745 86504 50773
rect 86344 50728 86504 50745
rect 101704 50959 101864 50976
rect 101704 50931 101739 50959
rect 101767 50931 101801 50959
rect 101829 50931 101864 50959
rect 101704 50897 101864 50931
rect 101704 50869 101739 50897
rect 101767 50869 101801 50897
rect 101829 50869 101864 50897
rect 101704 50835 101864 50869
rect 101704 50807 101739 50835
rect 101767 50807 101801 50835
rect 101829 50807 101864 50835
rect 101704 50773 101864 50807
rect 101704 50745 101739 50773
rect 101767 50745 101801 50773
rect 101829 50745 101864 50773
rect 101704 50728 101864 50745
rect 117064 50959 117224 50976
rect 117064 50931 117099 50959
rect 117127 50931 117161 50959
rect 117189 50931 117224 50959
rect 117064 50897 117224 50931
rect 117064 50869 117099 50897
rect 117127 50869 117161 50897
rect 117189 50869 117224 50897
rect 117064 50835 117224 50869
rect 117064 50807 117099 50835
rect 117127 50807 117161 50835
rect 117189 50807 117224 50835
rect 117064 50773 117224 50807
rect 117064 50745 117099 50773
rect 117127 50745 117161 50773
rect 117189 50745 117224 50773
rect 117064 50728 117224 50745
rect 132424 50959 132584 50976
rect 132424 50931 132459 50959
rect 132487 50931 132521 50959
rect 132549 50931 132584 50959
rect 132424 50897 132584 50931
rect 132424 50869 132459 50897
rect 132487 50869 132521 50897
rect 132549 50869 132584 50897
rect 132424 50835 132584 50869
rect 132424 50807 132459 50835
rect 132487 50807 132521 50835
rect 132549 50807 132584 50835
rect 132424 50773 132584 50807
rect 132424 50745 132459 50773
rect 132487 50745 132521 50773
rect 132549 50745 132584 50773
rect 132424 50728 132584 50745
rect 147784 50959 147944 50976
rect 147784 50931 147819 50959
rect 147847 50931 147881 50959
rect 147909 50931 147944 50959
rect 147784 50897 147944 50931
rect 147784 50869 147819 50897
rect 147847 50869 147881 50897
rect 147909 50869 147944 50897
rect 147784 50835 147944 50869
rect 147784 50807 147819 50835
rect 147847 50807 147881 50835
rect 147909 50807 147944 50835
rect 147784 50773 147944 50807
rect 147784 50745 147819 50773
rect 147847 50745 147881 50773
rect 147909 50745 147944 50773
rect 147784 50728 147944 50745
rect 163144 50959 163304 50976
rect 163144 50931 163179 50959
rect 163207 50931 163241 50959
rect 163269 50931 163304 50959
rect 163144 50897 163304 50931
rect 163144 50869 163179 50897
rect 163207 50869 163241 50897
rect 163269 50869 163304 50897
rect 163144 50835 163304 50869
rect 163144 50807 163179 50835
rect 163207 50807 163241 50835
rect 163269 50807 163304 50835
rect 163144 50773 163304 50807
rect 163144 50745 163179 50773
rect 163207 50745 163241 50773
rect 163269 50745 163304 50773
rect 163144 50728 163304 50745
rect 178504 50959 178664 50976
rect 178504 50931 178539 50959
rect 178567 50931 178601 50959
rect 178629 50931 178664 50959
rect 178504 50897 178664 50931
rect 178504 50869 178539 50897
rect 178567 50869 178601 50897
rect 178629 50869 178664 50897
rect 178504 50835 178664 50869
rect 178504 50807 178539 50835
rect 178567 50807 178601 50835
rect 178629 50807 178664 50835
rect 178504 50773 178664 50807
rect 178504 50745 178539 50773
rect 178567 50745 178601 50773
rect 178629 50745 178664 50773
rect 178504 50728 178664 50745
rect 193864 50959 194024 50976
rect 193864 50931 193899 50959
rect 193927 50931 193961 50959
rect 193989 50931 194024 50959
rect 193864 50897 194024 50931
rect 193864 50869 193899 50897
rect 193927 50869 193961 50897
rect 193989 50869 194024 50897
rect 193864 50835 194024 50869
rect 193864 50807 193899 50835
rect 193927 50807 193961 50835
rect 193989 50807 194024 50835
rect 193864 50773 194024 50807
rect 193864 50745 193899 50773
rect 193927 50745 193961 50773
rect 193989 50745 194024 50773
rect 193864 50728 194024 50745
rect 209224 50959 209384 50976
rect 209224 50931 209259 50959
rect 209287 50931 209321 50959
rect 209349 50931 209384 50959
rect 209224 50897 209384 50931
rect 209224 50869 209259 50897
rect 209287 50869 209321 50897
rect 209349 50869 209384 50897
rect 209224 50835 209384 50869
rect 209224 50807 209259 50835
rect 209287 50807 209321 50835
rect 209349 50807 209384 50835
rect 209224 50773 209384 50807
rect 209224 50745 209259 50773
rect 209287 50745 209321 50773
rect 209349 50745 209384 50773
rect 209224 50728 209384 50745
rect 224584 50959 224744 50976
rect 224584 50931 224619 50959
rect 224647 50931 224681 50959
rect 224709 50931 224744 50959
rect 224584 50897 224744 50931
rect 224584 50869 224619 50897
rect 224647 50869 224681 50897
rect 224709 50869 224744 50897
rect 224584 50835 224744 50869
rect 224584 50807 224619 50835
rect 224647 50807 224681 50835
rect 224709 50807 224744 50835
rect 224584 50773 224744 50807
rect 224584 50745 224619 50773
rect 224647 50745 224681 50773
rect 224709 50745 224744 50773
rect 224584 50728 224744 50745
rect 239944 50959 240104 50976
rect 239944 50931 239979 50959
rect 240007 50931 240041 50959
rect 240069 50931 240104 50959
rect 239944 50897 240104 50931
rect 239944 50869 239979 50897
rect 240007 50869 240041 50897
rect 240069 50869 240104 50897
rect 239944 50835 240104 50869
rect 239944 50807 239979 50835
rect 240007 50807 240041 50835
rect 240069 50807 240104 50835
rect 239944 50773 240104 50807
rect 239944 50745 239979 50773
rect 240007 50745 240041 50773
rect 240069 50745 240104 50773
rect 239944 50728 240104 50745
rect 32584 47959 32744 47976
rect 32584 47931 32619 47959
rect 32647 47931 32681 47959
rect 32709 47931 32744 47959
rect 32584 47897 32744 47931
rect 32584 47869 32619 47897
rect 32647 47869 32681 47897
rect 32709 47869 32744 47897
rect 32584 47835 32744 47869
rect 32584 47807 32619 47835
rect 32647 47807 32681 47835
rect 32709 47807 32744 47835
rect 32584 47773 32744 47807
rect 32584 47745 32619 47773
rect 32647 47745 32681 47773
rect 32709 47745 32744 47773
rect 32584 47728 32744 47745
rect 47944 47959 48104 47976
rect 47944 47931 47979 47959
rect 48007 47931 48041 47959
rect 48069 47931 48104 47959
rect 47944 47897 48104 47931
rect 47944 47869 47979 47897
rect 48007 47869 48041 47897
rect 48069 47869 48104 47897
rect 47944 47835 48104 47869
rect 47944 47807 47979 47835
rect 48007 47807 48041 47835
rect 48069 47807 48104 47835
rect 47944 47773 48104 47807
rect 47944 47745 47979 47773
rect 48007 47745 48041 47773
rect 48069 47745 48104 47773
rect 47944 47728 48104 47745
rect 63304 47959 63464 47976
rect 63304 47931 63339 47959
rect 63367 47931 63401 47959
rect 63429 47931 63464 47959
rect 63304 47897 63464 47931
rect 63304 47869 63339 47897
rect 63367 47869 63401 47897
rect 63429 47869 63464 47897
rect 63304 47835 63464 47869
rect 63304 47807 63339 47835
rect 63367 47807 63401 47835
rect 63429 47807 63464 47835
rect 63304 47773 63464 47807
rect 63304 47745 63339 47773
rect 63367 47745 63401 47773
rect 63429 47745 63464 47773
rect 63304 47728 63464 47745
rect 78664 47959 78824 47976
rect 78664 47931 78699 47959
rect 78727 47931 78761 47959
rect 78789 47931 78824 47959
rect 78664 47897 78824 47931
rect 78664 47869 78699 47897
rect 78727 47869 78761 47897
rect 78789 47869 78824 47897
rect 78664 47835 78824 47869
rect 78664 47807 78699 47835
rect 78727 47807 78761 47835
rect 78789 47807 78824 47835
rect 78664 47773 78824 47807
rect 78664 47745 78699 47773
rect 78727 47745 78761 47773
rect 78789 47745 78824 47773
rect 78664 47728 78824 47745
rect 94024 47959 94184 47976
rect 94024 47931 94059 47959
rect 94087 47931 94121 47959
rect 94149 47931 94184 47959
rect 94024 47897 94184 47931
rect 94024 47869 94059 47897
rect 94087 47869 94121 47897
rect 94149 47869 94184 47897
rect 94024 47835 94184 47869
rect 94024 47807 94059 47835
rect 94087 47807 94121 47835
rect 94149 47807 94184 47835
rect 94024 47773 94184 47807
rect 94024 47745 94059 47773
rect 94087 47745 94121 47773
rect 94149 47745 94184 47773
rect 94024 47728 94184 47745
rect 109384 47959 109544 47976
rect 109384 47931 109419 47959
rect 109447 47931 109481 47959
rect 109509 47931 109544 47959
rect 109384 47897 109544 47931
rect 109384 47869 109419 47897
rect 109447 47869 109481 47897
rect 109509 47869 109544 47897
rect 109384 47835 109544 47869
rect 109384 47807 109419 47835
rect 109447 47807 109481 47835
rect 109509 47807 109544 47835
rect 109384 47773 109544 47807
rect 109384 47745 109419 47773
rect 109447 47745 109481 47773
rect 109509 47745 109544 47773
rect 109384 47728 109544 47745
rect 124744 47959 124904 47976
rect 124744 47931 124779 47959
rect 124807 47931 124841 47959
rect 124869 47931 124904 47959
rect 124744 47897 124904 47931
rect 124744 47869 124779 47897
rect 124807 47869 124841 47897
rect 124869 47869 124904 47897
rect 124744 47835 124904 47869
rect 124744 47807 124779 47835
rect 124807 47807 124841 47835
rect 124869 47807 124904 47835
rect 124744 47773 124904 47807
rect 124744 47745 124779 47773
rect 124807 47745 124841 47773
rect 124869 47745 124904 47773
rect 124744 47728 124904 47745
rect 140104 47959 140264 47976
rect 140104 47931 140139 47959
rect 140167 47931 140201 47959
rect 140229 47931 140264 47959
rect 140104 47897 140264 47931
rect 140104 47869 140139 47897
rect 140167 47869 140201 47897
rect 140229 47869 140264 47897
rect 140104 47835 140264 47869
rect 140104 47807 140139 47835
rect 140167 47807 140201 47835
rect 140229 47807 140264 47835
rect 140104 47773 140264 47807
rect 140104 47745 140139 47773
rect 140167 47745 140201 47773
rect 140229 47745 140264 47773
rect 140104 47728 140264 47745
rect 155464 47959 155624 47976
rect 155464 47931 155499 47959
rect 155527 47931 155561 47959
rect 155589 47931 155624 47959
rect 155464 47897 155624 47931
rect 155464 47869 155499 47897
rect 155527 47869 155561 47897
rect 155589 47869 155624 47897
rect 155464 47835 155624 47869
rect 155464 47807 155499 47835
rect 155527 47807 155561 47835
rect 155589 47807 155624 47835
rect 155464 47773 155624 47807
rect 155464 47745 155499 47773
rect 155527 47745 155561 47773
rect 155589 47745 155624 47773
rect 155464 47728 155624 47745
rect 170824 47959 170984 47976
rect 170824 47931 170859 47959
rect 170887 47931 170921 47959
rect 170949 47931 170984 47959
rect 170824 47897 170984 47931
rect 170824 47869 170859 47897
rect 170887 47869 170921 47897
rect 170949 47869 170984 47897
rect 170824 47835 170984 47869
rect 170824 47807 170859 47835
rect 170887 47807 170921 47835
rect 170949 47807 170984 47835
rect 170824 47773 170984 47807
rect 170824 47745 170859 47773
rect 170887 47745 170921 47773
rect 170949 47745 170984 47773
rect 170824 47728 170984 47745
rect 186184 47959 186344 47976
rect 186184 47931 186219 47959
rect 186247 47931 186281 47959
rect 186309 47931 186344 47959
rect 186184 47897 186344 47931
rect 186184 47869 186219 47897
rect 186247 47869 186281 47897
rect 186309 47869 186344 47897
rect 186184 47835 186344 47869
rect 186184 47807 186219 47835
rect 186247 47807 186281 47835
rect 186309 47807 186344 47835
rect 186184 47773 186344 47807
rect 186184 47745 186219 47773
rect 186247 47745 186281 47773
rect 186309 47745 186344 47773
rect 186184 47728 186344 47745
rect 201544 47959 201704 47976
rect 201544 47931 201579 47959
rect 201607 47931 201641 47959
rect 201669 47931 201704 47959
rect 201544 47897 201704 47931
rect 201544 47869 201579 47897
rect 201607 47869 201641 47897
rect 201669 47869 201704 47897
rect 201544 47835 201704 47869
rect 201544 47807 201579 47835
rect 201607 47807 201641 47835
rect 201669 47807 201704 47835
rect 201544 47773 201704 47807
rect 201544 47745 201579 47773
rect 201607 47745 201641 47773
rect 201669 47745 201704 47773
rect 201544 47728 201704 47745
rect 216904 47959 217064 47976
rect 216904 47931 216939 47959
rect 216967 47931 217001 47959
rect 217029 47931 217064 47959
rect 216904 47897 217064 47931
rect 216904 47869 216939 47897
rect 216967 47869 217001 47897
rect 217029 47869 217064 47897
rect 216904 47835 217064 47869
rect 216904 47807 216939 47835
rect 216967 47807 217001 47835
rect 217029 47807 217064 47835
rect 216904 47773 217064 47807
rect 216904 47745 216939 47773
rect 216967 47745 217001 47773
rect 217029 47745 217064 47773
rect 216904 47728 217064 47745
rect 232264 47959 232424 47976
rect 232264 47931 232299 47959
rect 232327 47931 232361 47959
rect 232389 47931 232424 47959
rect 232264 47897 232424 47931
rect 232264 47869 232299 47897
rect 232327 47869 232361 47897
rect 232389 47869 232424 47897
rect 232264 47835 232424 47869
rect 232264 47807 232299 47835
rect 232327 47807 232361 47835
rect 232389 47807 232424 47835
rect 232264 47773 232424 47807
rect 232264 47745 232299 47773
rect 232327 47745 232361 47773
rect 232389 47745 232424 47773
rect 232264 47728 232424 47745
rect 247624 47959 247784 47976
rect 247624 47931 247659 47959
rect 247687 47931 247721 47959
rect 247749 47931 247784 47959
rect 247624 47897 247784 47931
rect 247624 47869 247659 47897
rect 247687 47869 247721 47897
rect 247749 47869 247784 47897
rect 247624 47835 247784 47869
rect 247624 47807 247659 47835
rect 247687 47807 247721 47835
rect 247749 47807 247784 47835
rect 247624 47773 247784 47807
rect 247624 47745 247659 47773
rect 247687 47745 247721 47773
rect 247749 47745 247784 47773
rect 247624 47728 247784 47745
rect 254529 47959 254839 56745
rect 254529 47931 254577 47959
rect 254605 47931 254639 47959
rect 254667 47931 254701 47959
rect 254729 47931 254763 47959
rect 254791 47931 254839 47959
rect 254529 47897 254839 47931
rect 254529 47869 254577 47897
rect 254605 47869 254639 47897
rect 254667 47869 254701 47897
rect 254729 47869 254763 47897
rect 254791 47869 254839 47897
rect 254529 47835 254839 47869
rect 254529 47807 254577 47835
rect 254605 47807 254639 47835
rect 254667 47807 254701 47835
rect 254729 47807 254763 47835
rect 254791 47807 254839 47835
rect 254529 47773 254839 47807
rect 254529 47745 254577 47773
rect 254605 47745 254639 47773
rect 254667 47745 254701 47773
rect 254729 47745 254763 47773
rect 254791 47745 254839 47773
rect 31389 41931 31437 41959
rect 31465 41931 31499 41959
rect 31527 41931 31561 41959
rect 31589 41931 31623 41959
rect 31651 41931 31699 41959
rect 31389 41897 31699 41931
rect 31389 41869 31437 41897
rect 31465 41869 31499 41897
rect 31527 41869 31561 41897
rect 31589 41869 31623 41897
rect 31651 41869 31699 41897
rect 31389 41835 31699 41869
rect 31389 41807 31437 41835
rect 31465 41807 31499 41835
rect 31527 41807 31561 41835
rect 31589 41807 31623 41835
rect 31651 41807 31699 41835
rect 31389 41773 31699 41807
rect 31389 41745 31437 41773
rect 31465 41745 31499 41773
rect 31527 41745 31561 41773
rect 31589 41745 31623 41773
rect 31651 41745 31699 41773
rect 31389 32959 31699 41745
rect 40264 41959 40424 41976
rect 40264 41931 40299 41959
rect 40327 41931 40361 41959
rect 40389 41931 40424 41959
rect 40264 41897 40424 41931
rect 40264 41869 40299 41897
rect 40327 41869 40361 41897
rect 40389 41869 40424 41897
rect 40264 41835 40424 41869
rect 40264 41807 40299 41835
rect 40327 41807 40361 41835
rect 40389 41807 40424 41835
rect 40264 41773 40424 41807
rect 40264 41745 40299 41773
rect 40327 41745 40361 41773
rect 40389 41745 40424 41773
rect 40264 41728 40424 41745
rect 55624 41959 55784 41976
rect 55624 41931 55659 41959
rect 55687 41931 55721 41959
rect 55749 41931 55784 41959
rect 55624 41897 55784 41931
rect 55624 41869 55659 41897
rect 55687 41869 55721 41897
rect 55749 41869 55784 41897
rect 55624 41835 55784 41869
rect 55624 41807 55659 41835
rect 55687 41807 55721 41835
rect 55749 41807 55784 41835
rect 55624 41773 55784 41807
rect 55624 41745 55659 41773
rect 55687 41745 55721 41773
rect 55749 41745 55784 41773
rect 55624 41728 55784 41745
rect 70984 41959 71144 41976
rect 70984 41931 71019 41959
rect 71047 41931 71081 41959
rect 71109 41931 71144 41959
rect 70984 41897 71144 41931
rect 70984 41869 71019 41897
rect 71047 41869 71081 41897
rect 71109 41869 71144 41897
rect 70984 41835 71144 41869
rect 70984 41807 71019 41835
rect 71047 41807 71081 41835
rect 71109 41807 71144 41835
rect 70984 41773 71144 41807
rect 70984 41745 71019 41773
rect 71047 41745 71081 41773
rect 71109 41745 71144 41773
rect 70984 41728 71144 41745
rect 86344 41959 86504 41976
rect 86344 41931 86379 41959
rect 86407 41931 86441 41959
rect 86469 41931 86504 41959
rect 86344 41897 86504 41931
rect 86344 41869 86379 41897
rect 86407 41869 86441 41897
rect 86469 41869 86504 41897
rect 86344 41835 86504 41869
rect 86344 41807 86379 41835
rect 86407 41807 86441 41835
rect 86469 41807 86504 41835
rect 86344 41773 86504 41807
rect 86344 41745 86379 41773
rect 86407 41745 86441 41773
rect 86469 41745 86504 41773
rect 86344 41728 86504 41745
rect 101704 41959 101864 41976
rect 101704 41931 101739 41959
rect 101767 41931 101801 41959
rect 101829 41931 101864 41959
rect 101704 41897 101864 41931
rect 101704 41869 101739 41897
rect 101767 41869 101801 41897
rect 101829 41869 101864 41897
rect 101704 41835 101864 41869
rect 101704 41807 101739 41835
rect 101767 41807 101801 41835
rect 101829 41807 101864 41835
rect 101704 41773 101864 41807
rect 101704 41745 101739 41773
rect 101767 41745 101801 41773
rect 101829 41745 101864 41773
rect 101704 41728 101864 41745
rect 117064 41959 117224 41976
rect 117064 41931 117099 41959
rect 117127 41931 117161 41959
rect 117189 41931 117224 41959
rect 117064 41897 117224 41931
rect 117064 41869 117099 41897
rect 117127 41869 117161 41897
rect 117189 41869 117224 41897
rect 117064 41835 117224 41869
rect 117064 41807 117099 41835
rect 117127 41807 117161 41835
rect 117189 41807 117224 41835
rect 117064 41773 117224 41807
rect 117064 41745 117099 41773
rect 117127 41745 117161 41773
rect 117189 41745 117224 41773
rect 117064 41728 117224 41745
rect 132424 41959 132584 41976
rect 132424 41931 132459 41959
rect 132487 41931 132521 41959
rect 132549 41931 132584 41959
rect 132424 41897 132584 41931
rect 132424 41869 132459 41897
rect 132487 41869 132521 41897
rect 132549 41869 132584 41897
rect 132424 41835 132584 41869
rect 132424 41807 132459 41835
rect 132487 41807 132521 41835
rect 132549 41807 132584 41835
rect 132424 41773 132584 41807
rect 132424 41745 132459 41773
rect 132487 41745 132521 41773
rect 132549 41745 132584 41773
rect 132424 41728 132584 41745
rect 147784 41959 147944 41976
rect 147784 41931 147819 41959
rect 147847 41931 147881 41959
rect 147909 41931 147944 41959
rect 147784 41897 147944 41931
rect 147784 41869 147819 41897
rect 147847 41869 147881 41897
rect 147909 41869 147944 41897
rect 147784 41835 147944 41869
rect 147784 41807 147819 41835
rect 147847 41807 147881 41835
rect 147909 41807 147944 41835
rect 147784 41773 147944 41807
rect 147784 41745 147819 41773
rect 147847 41745 147881 41773
rect 147909 41745 147944 41773
rect 147784 41728 147944 41745
rect 163144 41959 163304 41976
rect 163144 41931 163179 41959
rect 163207 41931 163241 41959
rect 163269 41931 163304 41959
rect 163144 41897 163304 41931
rect 163144 41869 163179 41897
rect 163207 41869 163241 41897
rect 163269 41869 163304 41897
rect 163144 41835 163304 41869
rect 163144 41807 163179 41835
rect 163207 41807 163241 41835
rect 163269 41807 163304 41835
rect 163144 41773 163304 41807
rect 163144 41745 163179 41773
rect 163207 41745 163241 41773
rect 163269 41745 163304 41773
rect 163144 41728 163304 41745
rect 178504 41959 178664 41976
rect 178504 41931 178539 41959
rect 178567 41931 178601 41959
rect 178629 41931 178664 41959
rect 178504 41897 178664 41931
rect 178504 41869 178539 41897
rect 178567 41869 178601 41897
rect 178629 41869 178664 41897
rect 178504 41835 178664 41869
rect 178504 41807 178539 41835
rect 178567 41807 178601 41835
rect 178629 41807 178664 41835
rect 178504 41773 178664 41807
rect 178504 41745 178539 41773
rect 178567 41745 178601 41773
rect 178629 41745 178664 41773
rect 178504 41728 178664 41745
rect 193864 41959 194024 41976
rect 193864 41931 193899 41959
rect 193927 41931 193961 41959
rect 193989 41931 194024 41959
rect 193864 41897 194024 41931
rect 193864 41869 193899 41897
rect 193927 41869 193961 41897
rect 193989 41869 194024 41897
rect 193864 41835 194024 41869
rect 193864 41807 193899 41835
rect 193927 41807 193961 41835
rect 193989 41807 194024 41835
rect 193864 41773 194024 41807
rect 193864 41745 193899 41773
rect 193927 41745 193961 41773
rect 193989 41745 194024 41773
rect 193864 41728 194024 41745
rect 209224 41959 209384 41976
rect 209224 41931 209259 41959
rect 209287 41931 209321 41959
rect 209349 41931 209384 41959
rect 209224 41897 209384 41931
rect 209224 41869 209259 41897
rect 209287 41869 209321 41897
rect 209349 41869 209384 41897
rect 209224 41835 209384 41869
rect 209224 41807 209259 41835
rect 209287 41807 209321 41835
rect 209349 41807 209384 41835
rect 209224 41773 209384 41807
rect 209224 41745 209259 41773
rect 209287 41745 209321 41773
rect 209349 41745 209384 41773
rect 209224 41728 209384 41745
rect 224584 41959 224744 41976
rect 224584 41931 224619 41959
rect 224647 41931 224681 41959
rect 224709 41931 224744 41959
rect 224584 41897 224744 41931
rect 224584 41869 224619 41897
rect 224647 41869 224681 41897
rect 224709 41869 224744 41897
rect 224584 41835 224744 41869
rect 224584 41807 224619 41835
rect 224647 41807 224681 41835
rect 224709 41807 224744 41835
rect 224584 41773 224744 41807
rect 224584 41745 224619 41773
rect 224647 41745 224681 41773
rect 224709 41745 224744 41773
rect 224584 41728 224744 41745
rect 239944 41959 240104 41976
rect 239944 41931 239979 41959
rect 240007 41931 240041 41959
rect 240069 41931 240104 41959
rect 239944 41897 240104 41931
rect 239944 41869 239979 41897
rect 240007 41869 240041 41897
rect 240069 41869 240104 41897
rect 239944 41835 240104 41869
rect 239944 41807 239979 41835
rect 240007 41807 240041 41835
rect 240069 41807 240104 41835
rect 239944 41773 240104 41807
rect 239944 41745 239979 41773
rect 240007 41745 240041 41773
rect 240069 41745 240104 41773
rect 239944 41728 240104 41745
rect 32584 38959 32744 38976
rect 32584 38931 32619 38959
rect 32647 38931 32681 38959
rect 32709 38931 32744 38959
rect 32584 38897 32744 38931
rect 32584 38869 32619 38897
rect 32647 38869 32681 38897
rect 32709 38869 32744 38897
rect 32584 38835 32744 38869
rect 32584 38807 32619 38835
rect 32647 38807 32681 38835
rect 32709 38807 32744 38835
rect 32584 38773 32744 38807
rect 32584 38745 32619 38773
rect 32647 38745 32681 38773
rect 32709 38745 32744 38773
rect 32584 38728 32744 38745
rect 47944 38959 48104 38976
rect 47944 38931 47979 38959
rect 48007 38931 48041 38959
rect 48069 38931 48104 38959
rect 47944 38897 48104 38931
rect 47944 38869 47979 38897
rect 48007 38869 48041 38897
rect 48069 38869 48104 38897
rect 47944 38835 48104 38869
rect 47944 38807 47979 38835
rect 48007 38807 48041 38835
rect 48069 38807 48104 38835
rect 47944 38773 48104 38807
rect 47944 38745 47979 38773
rect 48007 38745 48041 38773
rect 48069 38745 48104 38773
rect 47944 38728 48104 38745
rect 63304 38959 63464 38976
rect 63304 38931 63339 38959
rect 63367 38931 63401 38959
rect 63429 38931 63464 38959
rect 63304 38897 63464 38931
rect 63304 38869 63339 38897
rect 63367 38869 63401 38897
rect 63429 38869 63464 38897
rect 63304 38835 63464 38869
rect 63304 38807 63339 38835
rect 63367 38807 63401 38835
rect 63429 38807 63464 38835
rect 63304 38773 63464 38807
rect 63304 38745 63339 38773
rect 63367 38745 63401 38773
rect 63429 38745 63464 38773
rect 63304 38728 63464 38745
rect 78664 38959 78824 38976
rect 78664 38931 78699 38959
rect 78727 38931 78761 38959
rect 78789 38931 78824 38959
rect 78664 38897 78824 38931
rect 78664 38869 78699 38897
rect 78727 38869 78761 38897
rect 78789 38869 78824 38897
rect 78664 38835 78824 38869
rect 78664 38807 78699 38835
rect 78727 38807 78761 38835
rect 78789 38807 78824 38835
rect 78664 38773 78824 38807
rect 78664 38745 78699 38773
rect 78727 38745 78761 38773
rect 78789 38745 78824 38773
rect 78664 38728 78824 38745
rect 94024 38959 94184 38976
rect 94024 38931 94059 38959
rect 94087 38931 94121 38959
rect 94149 38931 94184 38959
rect 94024 38897 94184 38931
rect 94024 38869 94059 38897
rect 94087 38869 94121 38897
rect 94149 38869 94184 38897
rect 94024 38835 94184 38869
rect 94024 38807 94059 38835
rect 94087 38807 94121 38835
rect 94149 38807 94184 38835
rect 94024 38773 94184 38807
rect 94024 38745 94059 38773
rect 94087 38745 94121 38773
rect 94149 38745 94184 38773
rect 94024 38728 94184 38745
rect 109384 38959 109544 38976
rect 109384 38931 109419 38959
rect 109447 38931 109481 38959
rect 109509 38931 109544 38959
rect 109384 38897 109544 38931
rect 109384 38869 109419 38897
rect 109447 38869 109481 38897
rect 109509 38869 109544 38897
rect 109384 38835 109544 38869
rect 109384 38807 109419 38835
rect 109447 38807 109481 38835
rect 109509 38807 109544 38835
rect 109384 38773 109544 38807
rect 109384 38745 109419 38773
rect 109447 38745 109481 38773
rect 109509 38745 109544 38773
rect 109384 38728 109544 38745
rect 124744 38959 124904 38976
rect 124744 38931 124779 38959
rect 124807 38931 124841 38959
rect 124869 38931 124904 38959
rect 124744 38897 124904 38931
rect 124744 38869 124779 38897
rect 124807 38869 124841 38897
rect 124869 38869 124904 38897
rect 124744 38835 124904 38869
rect 124744 38807 124779 38835
rect 124807 38807 124841 38835
rect 124869 38807 124904 38835
rect 124744 38773 124904 38807
rect 124744 38745 124779 38773
rect 124807 38745 124841 38773
rect 124869 38745 124904 38773
rect 124744 38728 124904 38745
rect 140104 38959 140264 38976
rect 140104 38931 140139 38959
rect 140167 38931 140201 38959
rect 140229 38931 140264 38959
rect 140104 38897 140264 38931
rect 140104 38869 140139 38897
rect 140167 38869 140201 38897
rect 140229 38869 140264 38897
rect 140104 38835 140264 38869
rect 140104 38807 140139 38835
rect 140167 38807 140201 38835
rect 140229 38807 140264 38835
rect 140104 38773 140264 38807
rect 140104 38745 140139 38773
rect 140167 38745 140201 38773
rect 140229 38745 140264 38773
rect 140104 38728 140264 38745
rect 155464 38959 155624 38976
rect 155464 38931 155499 38959
rect 155527 38931 155561 38959
rect 155589 38931 155624 38959
rect 155464 38897 155624 38931
rect 155464 38869 155499 38897
rect 155527 38869 155561 38897
rect 155589 38869 155624 38897
rect 155464 38835 155624 38869
rect 155464 38807 155499 38835
rect 155527 38807 155561 38835
rect 155589 38807 155624 38835
rect 155464 38773 155624 38807
rect 155464 38745 155499 38773
rect 155527 38745 155561 38773
rect 155589 38745 155624 38773
rect 155464 38728 155624 38745
rect 170824 38959 170984 38976
rect 170824 38931 170859 38959
rect 170887 38931 170921 38959
rect 170949 38931 170984 38959
rect 170824 38897 170984 38931
rect 170824 38869 170859 38897
rect 170887 38869 170921 38897
rect 170949 38869 170984 38897
rect 170824 38835 170984 38869
rect 170824 38807 170859 38835
rect 170887 38807 170921 38835
rect 170949 38807 170984 38835
rect 170824 38773 170984 38807
rect 170824 38745 170859 38773
rect 170887 38745 170921 38773
rect 170949 38745 170984 38773
rect 170824 38728 170984 38745
rect 186184 38959 186344 38976
rect 186184 38931 186219 38959
rect 186247 38931 186281 38959
rect 186309 38931 186344 38959
rect 186184 38897 186344 38931
rect 186184 38869 186219 38897
rect 186247 38869 186281 38897
rect 186309 38869 186344 38897
rect 186184 38835 186344 38869
rect 186184 38807 186219 38835
rect 186247 38807 186281 38835
rect 186309 38807 186344 38835
rect 186184 38773 186344 38807
rect 186184 38745 186219 38773
rect 186247 38745 186281 38773
rect 186309 38745 186344 38773
rect 186184 38728 186344 38745
rect 201544 38959 201704 38976
rect 201544 38931 201579 38959
rect 201607 38931 201641 38959
rect 201669 38931 201704 38959
rect 201544 38897 201704 38931
rect 201544 38869 201579 38897
rect 201607 38869 201641 38897
rect 201669 38869 201704 38897
rect 201544 38835 201704 38869
rect 201544 38807 201579 38835
rect 201607 38807 201641 38835
rect 201669 38807 201704 38835
rect 201544 38773 201704 38807
rect 201544 38745 201579 38773
rect 201607 38745 201641 38773
rect 201669 38745 201704 38773
rect 201544 38728 201704 38745
rect 216904 38959 217064 38976
rect 216904 38931 216939 38959
rect 216967 38931 217001 38959
rect 217029 38931 217064 38959
rect 216904 38897 217064 38931
rect 216904 38869 216939 38897
rect 216967 38869 217001 38897
rect 217029 38869 217064 38897
rect 216904 38835 217064 38869
rect 216904 38807 216939 38835
rect 216967 38807 217001 38835
rect 217029 38807 217064 38835
rect 216904 38773 217064 38807
rect 216904 38745 216939 38773
rect 216967 38745 217001 38773
rect 217029 38745 217064 38773
rect 216904 38728 217064 38745
rect 232264 38959 232424 38976
rect 232264 38931 232299 38959
rect 232327 38931 232361 38959
rect 232389 38931 232424 38959
rect 232264 38897 232424 38931
rect 232264 38869 232299 38897
rect 232327 38869 232361 38897
rect 232389 38869 232424 38897
rect 232264 38835 232424 38869
rect 232264 38807 232299 38835
rect 232327 38807 232361 38835
rect 232389 38807 232424 38835
rect 232264 38773 232424 38807
rect 232264 38745 232299 38773
rect 232327 38745 232361 38773
rect 232389 38745 232424 38773
rect 232264 38728 232424 38745
rect 247624 38959 247784 38976
rect 247624 38931 247659 38959
rect 247687 38931 247721 38959
rect 247749 38931 247784 38959
rect 247624 38897 247784 38931
rect 247624 38869 247659 38897
rect 247687 38869 247721 38897
rect 247749 38869 247784 38897
rect 247624 38835 247784 38869
rect 247624 38807 247659 38835
rect 247687 38807 247721 38835
rect 247749 38807 247784 38835
rect 247624 38773 247784 38807
rect 247624 38745 247659 38773
rect 247687 38745 247721 38773
rect 247749 38745 247784 38773
rect 247624 38728 247784 38745
rect 254529 38959 254839 47745
rect 254529 38931 254577 38959
rect 254605 38931 254639 38959
rect 254667 38931 254701 38959
rect 254729 38931 254763 38959
rect 254791 38931 254839 38959
rect 254529 38897 254839 38931
rect 254529 38869 254577 38897
rect 254605 38869 254639 38897
rect 254667 38869 254701 38897
rect 254729 38869 254763 38897
rect 254791 38869 254839 38897
rect 254529 38835 254839 38869
rect 254529 38807 254577 38835
rect 254605 38807 254639 38835
rect 254667 38807 254701 38835
rect 254729 38807 254763 38835
rect 254791 38807 254839 38835
rect 254529 38773 254839 38807
rect 254529 38745 254577 38773
rect 254605 38745 254639 38773
rect 254667 38745 254701 38773
rect 254729 38745 254763 38773
rect 254791 38745 254839 38773
rect 31389 32931 31437 32959
rect 31465 32931 31499 32959
rect 31527 32931 31561 32959
rect 31589 32931 31623 32959
rect 31651 32931 31699 32959
rect 31389 32897 31699 32931
rect 31389 32869 31437 32897
rect 31465 32869 31499 32897
rect 31527 32869 31561 32897
rect 31589 32869 31623 32897
rect 31651 32869 31699 32897
rect 31389 32835 31699 32869
rect 31389 32807 31437 32835
rect 31465 32807 31499 32835
rect 31527 32807 31561 32835
rect 31589 32807 31623 32835
rect 31651 32807 31699 32835
rect 31389 32773 31699 32807
rect 31389 32745 31437 32773
rect 31465 32745 31499 32773
rect 31527 32745 31561 32773
rect 31589 32745 31623 32773
rect 31651 32745 31699 32773
rect 31389 23959 31699 32745
rect 40264 32959 40424 32976
rect 40264 32931 40299 32959
rect 40327 32931 40361 32959
rect 40389 32931 40424 32959
rect 40264 32897 40424 32931
rect 40264 32869 40299 32897
rect 40327 32869 40361 32897
rect 40389 32869 40424 32897
rect 40264 32835 40424 32869
rect 40264 32807 40299 32835
rect 40327 32807 40361 32835
rect 40389 32807 40424 32835
rect 40264 32773 40424 32807
rect 40264 32745 40299 32773
rect 40327 32745 40361 32773
rect 40389 32745 40424 32773
rect 40264 32728 40424 32745
rect 55624 32959 55784 32976
rect 55624 32931 55659 32959
rect 55687 32931 55721 32959
rect 55749 32931 55784 32959
rect 55624 32897 55784 32931
rect 55624 32869 55659 32897
rect 55687 32869 55721 32897
rect 55749 32869 55784 32897
rect 55624 32835 55784 32869
rect 55624 32807 55659 32835
rect 55687 32807 55721 32835
rect 55749 32807 55784 32835
rect 55624 32773 55784 32807
rect 55624 32745 55659 32773
rect 55687 32745 55721 32773
rect 55749 32745 55784 32773
rect 55624 32728 55784 32745
rect 70984 32959 71144 32976
rect 70984 32931 71019 32959
rect 71047 32931 71081 32959
rect 71109 32931 71144 32959
rect 70984 32897 71144 32931
rect 70984 32869 71019 32897
rect 71047 32869 71081 32897
rect 71109 32869 71144 32897
rect 70984 32835 71144 32869
rect 70984 32807 71019 32835
rect 71047 32807 71081 32835
rect 71109 32807 71144 32835
rect 70984 32773 71144 32807
rect 70984 32745 71019 32773
rect 71047 32745 71081 32773
rect 71109 32745 71144 32773
rect 70984 32728 71144 32745
rect 86344 32959 86504 32976
rect 86344 32931 86379 32959
rect 86407 32931 86441 32959
rect 86469 32931 86504 32959
rect 86344 32897 86504 32931
rect 86344 32869 86379 32897
rect 86407 32869 86441 32897
rect 86469 32869 86504 32897
rect 86344 32835 86504 32869
rect 86344 32807 86379 32835
rect 86407 32807 86441 32835
rect 86469 32807 86504 32835
rect 86344 32773 86504 32807
rect 86344 32745 86379 32773
rect 86407 32745 86441 32773
rect 86469 32745 86504 32773
rect 86344 32728 86504 32745
rect 101704 32959 101864 32976
rect 101704 32931 101739 32959
rect 101767 32931 101801 32959
rect 101829 32931 101864 32959
rect 101704 32897 101864 32931
rect 101704 32869 101739 32897
rect 101767 32869 101801 32897
rect 101829 32869 101864 32897
rect 101704 32835 101864 32869
rect 101704 32807 101739 32835
rect 101767 32807 101801 32835
rect 101829 32807 101864 32835
rect 101704 32773 101864 32807
rect 101704 32745 101739 32773
rect 101767 32745 101801 32773
rect 101829 32745 101864 32773
rect 101704 32728 101864 32745
rect 117064 32959 117224 32976
rect 117064 32931 117099 32959
rect 117127 32931 117161 32959
rect 117189 32931 117224 32959
rect 117064 32897 117224 32931
rect 117064 32869 117099 32897
rect 117127 32869 117161 32897
rect 117189 32869 117224 32897
rect 117064 32835 117224 32869
rect 117064 32807 117099 32835
rect 117127 32807 117161 32835
rect 117189 32807 117224 32835
rect 117064 32773 117224 32807
rect 117064 32745 117099 32773
rect 117127 32745 117161 32773
rect 117189 32745 117224 32773
rect 117064 32728 117224 32745
rect 132424 32959 132584 32976
rect 132424 32931 132459 32959
rect 132487 32931 132521 32959
rect 132549 32931 132584 32959
rect 132424 32897 132584 32931
rect 132424 32869 132459 32897
rect 132487 32869 132521 32897
rect 132549 32869 132584 32897
rect 132424 32835 132584 32869
rect 132424 32807 132459 32835
rect 132487 32807 132521 32835
rect 132549 32807 132584 32835
rect 132424 32773 132584 32807
rect 132424 32745 132459 32773
rect 132487 32745 132521 32773
rect 132549 32745 132584 32773
rect 132424 32728 132584 32745
rect 147784 32959 147944 32976
rect 147784 32931 147819 32959
rect 147847 32931 147881 32959
rect 147909 32931 147944 32959
rect 147784 32897 147944 32931
rect 147784 32869 147819 32897
rect 147847 32869 147881 32897
rect 147909 32869 147944 32897
rect 147784 32835 147944 32869
rect 147784 32807 147819 32835
rect 147847 32807 147881 32835
rect 147909 32807 147944 32835
rect 147784 32773 147944 32807
rect 147784 32745 147819 32773
rect 147847 32745 147881 32773
rect 147909 32745 147944 32773
rect 147784 32728 147944 32745
rect 163144 32959 163304 32976
rect 163144 32931 163179 32959
rect 163207 32931 163241 32959
rect 163269 32931 163304 32959
rect 163144 32897 163304 32931
rect 163144 32869 163179 32897
rect 163207 32869 163241 32897
rect 163269 32869 163304 32897
rect 163144 32835 163304 32869
rect 163144 32807 163179 32835
rect 163207 32807 163241 32835
rect 163269 32807 163304 32835
rect 163144 32773 163304 32807
rect 163144 32745 163179 32773
rect 163207 32745 163241 32773
rect 163269 32745 163304 32773
rect 163144 32728 163304 32745
rect 178504 32959 178664 32976
rect 178504 32931 178539 32959
rect 178567 32931 178601 32959
rect 178629 32931 178664 32959
rect 178504 32897 178664 32931
rect 178504 32869 178539 32897
rect 178567 32869 178601 32897
rect 178629 32869 178664 32897
rect 178504 32835 178664 32869
rect 178504 32807 178539 32835
rect 178567 32807 178601 32835
rect 178629 32807 178664 32835
rect 178504 32773 178664 32807
rect 178504 32745 178539 32773
rect 178567 32745 178601 32773
rect 178629 32745 178664 32773
rect 178504 32728 178664 32745
rect 193864 32959 194024 32976
rect 193864 32931 193899 32959
rect 193927 32931 193961 32959
rect 193989 32931 194024 32959
rect 193864 32897 194024 32931
rect 193864 32869 193899 32897
rect 193927 32869 193961 32897
rect 193989 32869 194024 32897
rect 193864 32835 194024 32869
rect 193864 32807 193899 32835
rect 193927 32807 193961 32835
rect 193989 32807 194024 32835
rect 193864 32773 194024 32807
rect 193864 32745 193899 32773
rect 193927 32745 193961 32773
rect 193989 32745 194024 32773
rect 193864 32728 194024 32745
rect 209224 32959 209384 32976
rect 209224 32931 209259 32959
rect 209287 32931 209321 32959
rect 209349 32931 209384 32959
rect 209224 32897 209384 32931
rect 209224 32869 209259 32897
rect 209287 32869 209321 32897
rect 209349 32869 209384 32897
rect 209224 32835 209384 32869
rect 209224 32807 209259 32835
rect 209287 32807 209321 32835
rect 209349 32807 209384 32835
rect 209224 32773 209384 32807
rect 209224 32745 209259 32773
rect 209287 32745 209321 32773
rect 209349 32745 209384 32773
rect 209224 32728 209384 32745
rect 224584 32959 224744 32976
rect 224584 32931 224619 32959
rect 224647 32931 224681 32959
rect 224709 32931 224744 32959
rect 224584 32897 224744 32931
rect 224584 32869 224619 32897
rect 224647 32869 224681 32897
rect 224709 32869 224744 32897
rect 224584 32835 224744 32869
rect 224584 32807 224619 32835
rect 224647 32807 224681 32835
rect 224709 32807 224744 32835
rect 224584 32773 224744 32807
rect 224584 32745 224619 32773
rect 224647 32745 224681 32773
rect 224709 32745 224744 32773
rect 224584 32728 224744 32745
rect 239944 32959 240104 32976
rect 239944 32931 239979 32959
rect 240007 32931 240041 32959
rect 240069 32931 240104 32959
rect 239944 32897 240104 32931
rect 239944 32869 239979 32897
rect 240007 32869 240041 32897
rect 240069 32869 240104 32897
rect 239944 32835 240104 32869
rect 239944 32807 239979 32835
rect 240007 32807 240041 32835
rect 240069 32807 240104 32835
rect 239944 32773 240104 32807
rect 239944 32745 239979 32773
rect 240007 32745 240041 32773
rect 240069 32745 240104 32773
rect 239944 32728 240104 32745
rect 32584 29959 32744 29976
rect 32584 29931 32619 29959
rect 32647 29931 32681 29959
rect 32709 29931 32744 29959
rect 32584 29897 32744 29931
rect 32584 29869 32619 29897
rect 32647 29869 32681 29897
rect 32709 29869 32744 29897
rect 32584 29835 32744 29869
rect 32584 29807 32619 29835
rect 32647 29807 32681 29835
rect 32709 29807 32744 29835
rect 32584 29773 32744 29807
rect 32584 29745 32619 29773
rect 32647 29745 32681 29773
rect 32709 29745 32744 29773
rect 32584 29728 32744 29745
rect 47944 29959 48104 29976
rect 47944 29931 47979 29959
rect 48007 29931 48041 29959
rect 48069 29931 48104 29959
rect 47944 29897 48104 29931
rect 47944 29869 47979 29897
rect 48007 29869 48041 29897
rect 48069 29869 48104 29897
rect 47944 29835 48104 29869
rect 47944 29807 47979 29835
rect 48007 29807 48041 29835
rect 48069 29807 48104 29835
rect 47944 29773 48104 29807
rect 47944 29745 47979 29773
rect 48007 29745 48041 29773
rect 48069 29745 48104 29773
rect 47944 29728 48104 29745
rect 63304 29959 63464 29976
rect 63304 29931 63339 29959
rect 63367 29931 63401 29959
rect 63429 29931 63464 29959
rect 63304 29897 63464 29931
rect 63304 29869 63339 29897
rect 63367 29869 63401 29897
rect 63429 29869 63464 29897
rect 63304 29835 63464 29869
rect 63304 29807 63339 29835
rect 63367 29807 63401 29835
rect 63429 29807 63464 29835
rect 63304 29773 63464 29807
rect 63304 29745 63339 29773
rect 63367 29745 63401 29773
rect 63429 29745 63464 29773
rect 63304 29728 63464 29745
rect 78664 29959 78824 29976
rect 78664 29931 78699 29959
rect 78727 29931 78761 29959
rect 78789 29931 78824 29959
rect 78664 29897 78824 29931
rect 78664 29869 78699 29897
rect 78727 29869 78761 29897
rect 78789 29869 78824 29897
rect 78664 29835 78824 29869
rect 78664 29807 78699 29835
rect 78727 29807 78761 29835
rect 78789 29807 78824 29835
rect 78664 29773 78824 29807
rect 78664 29745 78699 29773
rect 78727 29745 78761 29773
rect 78789 29745 78824 29773
rect 78664 29728 78824 29745
rect 94024 29959 94184 29976
rect 94024 29931 94059 29959
rect 94087 29931 94121 29959
rect 94149 29931 94184 29959
rect 94024 29897 94184 29931
rect 94024 29869 94059 29897
rect 94087 29869 94121 29897
rect 94149 29869 94184 29897
rect 94024 29835 94184 29869
rect 94024 29807 94059 29835
rect 94087 29807 94121 29835
rect 94149 29807 94184 29835
rect 94024 29773 94184 29807
rect 94024 29745 94059 29773
rect 94087 29745 94121 29773
rect 94149 29745 94184 29773
rect 94024 29728 94184 29745
rect 109384 29959 109544 29976
rect 109384 29931 109419 29959
rect 109447 29931 109481 29959
rect 109509 29931 109544 29959
rect 109384 29897 109544 29931
rect 109384 29869 109419 29897
rect 109447 29869 109481 29897
rect 109509 29869 109544 29897
rect 109384 29835 109544 29869
rect 109384 29807 109419 29835
rect 109447 29807 109481 29835
rect 109509 29807 109544 29835
rect 109384 29773 109544 29807
rect 109384 29745 109419 29773
rect 109447 29745 109481 29773
rect 109509 29745 109544 29773
rect 109384 29728 109544 29745
rect 124744 29959 124904 29976
rect 124744 29931 124779 29959
rect 124807 29931 124841 29959
rect 124869 29931 124904 29959
rect 124744 29897 124904 29931
rect 124744 29869 124779 29897
rect 124807 29869 124841 29897
rect 124869 29869 124904 29897
rect 124744 29835 124904 29869
rect 124744 29807 124779 29835
rect 124807 29807 124841 29835
rect 124869 29807 124904 29835
rect 124744 29773 124904 29807
rect 124744 29745 124779 29773
rect 124807 29745 124841 29773
rect 124869 29745 124904 29773
rect 124744 29728 124904 29745
rect 140104 29959 140264 29976
rect 140104 29931 140139 29959
rect 140167 29931 140201 29959
rect 140229 29931 140264 29959
rect 140104 29897 140264 29931
rect 140104 29869 140139 29897
rect 140167 29869 140201 29897
rect 140229 29869 140264 29897
rect 140104 29835 140264 29869
rect 140104 29807 140139 29835
rect 140167 29807 140201 29835
rect 140229 29807 140264 29835
rect 140104 29773 140264 29807
rect 140104 29745 140139 29773
rect 140167 29745 140201 29773
rect 140229 29745 140264 29773
rect 140104 29728 140264 29745
rect 155464 29959 155624 29976
rect 155464 29931 155499 29959
rect 155527 29931 155561 29959
rect 155589 29931 155624 29959
rect 155464 29897 155624 29931
rect 155464 29869 155499 29897
rect 155527 29869 155561 29897
rect 155589 29869 155624 29897
rect 155464 29835 155624 29869
rect 155464 29807 155499 29835
rect 155527 29807 155561 29835
rect 155589 29807 155624 29835
rect 155464 29773 155624 29807
rect 155464 29745 155499 29773
rect 155527 29745 155561 29773
rect 155589 29745 155624 29773
rect 155464 29728 155624 29745
rect 170824 29959 170984 29976
rect 170824 29931 170859 29959
rect 170887 29931 170921 29959
rect 170949 29931 170984 29959
rect 170824 29897 170984 29931
rect 170824 29869 170859 29897
rect 170887 29869 170921 29897
rect 170949 29869 170984 29897
rect 170824 29835 170984 29869
rect 170824 29807 170859 29835
rect 170887 29807 170921 29835
rect 170949 29807 170984 29835
rect 170824 29773 170984 29807
rect 170824 29745 170859 29773
rect 170887 29745 170921 29773
rect 170949 29745 170984 29773
rect 170824 29728 170984 29745
rect 186184 29959 186344 29976
rect 186184 29931 186219 29959
rect 186247 29931 186281 29959
rect 186309 29931 186344 29959
rect 186184 29897 186344 29931
rect 186184 29869 186219 29897
rect 186247 29869 186281 29897
rect 186309 29869 186344 29897
rect 186184 29835 186344 29869
rect 186184 29807 186219 29835
rect 186247 29807 186281 29835
rect 186309 29807 186344 29835
rect 186184 29773 186344 29807
rect 186184 29745 186219 29773
rect 186247 29745 186281 29773
rect 186309 29745 186344 29773
rect 186184 29728 186344 29745
rect 201544 29959 201704 29976
rect 201544 29931 201579 29959
rect 201607 29931 201641 29959
rect 201669 29931 201704 29959
rect 201544 29897 201704 29931
rect 201544 29869 201579 29897
rect 201607 29869 201641 29897
rect 201669 29869 201704 29897
rect 201544 29835 201704 29869
rect 201544 29807 201579 29835
rect 201607 29807 201641 29835
rect 201669 29807 201704 29835
rect 201544 29773 201704 29807
rect 201544 29745 201579 29773
rect 201607 29745 201641 29773
rect 201669 29745 201704 29773
rect 201544 29728 201704 29745
rect 216904 29959 217064 29976
rect 216904 29931 216939 29959
rect 216967 29931 217001 29959
rect 217029 29931 217064 29959
rect 216904 29897 217064 29931
rect 216904 29869 216939 29897
rect 216967 29869 217001 29897
rect 217029 29869 217064 29897
rect 216904 29835 217064 29869
rect 216904 29807 216939 29835
rect 216967 29807 217001 29835
rect 217029 29807 217064 29835
rect 216904 29773 217064 29807
rect 216904 29745 216939 29773
rect 216967 29745 217001 29773
rect 217029 29745 217064 29773
rect 216904 29728 217064 29745
rect 232264 29959 232424 29976
rect 232264 29931 232299 29959
rect 232327 29931 232361 29959
rect 232389 29931 232424 29959
rect 232264 29897 232424 29931
rect 232264 29869 232299 29897
rect 232327 29869 232361 29897
rect 232389 29869 232424 29897
rect 232264 29835 232424 29869
rect 232264 29807 232299 29835
rect 232327 29807 232361 29835
rect 232389 29807 232424 29835
rect 232264 29773 232424 29807
rect 232264 29745 232299 29773
rect 232327 29745 232361 29773
rect 232389 29745 232424 29773
rect 232264 29728 232424 29745
rect 247624 29959 247784 29976
rect 247624 29931 247659 29959
rect 247687 29931 247721 29959
rect 247749 29931 247784 29959
rect 247624 29897 247784 29931
rect 247624 29869 247659 29897
rect 247687 29869 247721 29897
rect 247749 29869 247784 29897
rect 247624 29835 247784 29869
rect 247624 29807 247659 29835
rect 247687 29807 247721 29835
rect 247749 29807 247784 29835
rect 247624 29773 247784 29807
rect 247624 29745 247659 29773
rect 247687 29745 247721 29773
rect 247749 29745 247784 29773
rect 247624 29728 247784 29745
rect 254529 29959 254839 38745
rect 254529 29931 254577 29959
rect 254605 29931 254639 29959
rect 254667 29931 254701 29959
rect 254729 29931 254763 29959
rect 254791 29931 254839 29959
rect 254529 29897 254839 29931
rect 254529 29869 254577 29897
rect 254605 29869 254639 29897
rect 254667 29869 254701 29897
rect 254729 29869 254763 29897
rect 254791 29869 254839 29897
rect 254529 29835 254839 29869
rect 254529 29807 254577 29835
rect 254605 29807 254639 29835
rect 254667 29807 254701 29835
rect 254729 29807 254763 29835
rect 254791 29807 254839 29835
rect 254529 29773 254839 29807
rect 254529 29745 254577 29773
rect 254605 29745 254639 29773
rect 254667 29745 254701 29773
rect 254729 29745 254763 29773
rect 254791 29745 254839 29773
rect 31389 23931 31437 23959
rect 31465 23931 31499 23959
rect 31527 23931 31561 23959
rect 31589 23931 31623 23959
rect 31651 23931 31699 23959
rect 31389 23897 31699 23931
rect 31389 23869 31437 23897
rect 31465 23869 31499 23897
rect 31527 23869 31561 23897
rect 31589 23869 31623 23897
rect 31651 23869 31699 23897
rect 31389 23835 31699 23869
rect 31389 23807 31437 23835
rect 31465 23807 31499 23835
rect 31527 23807 31561 23835
rect 31589 23807 31623 23835
rect 31651 23807 31699 23835
rect 31389 23773 31699 23807
rect 31389 23745 31437 23773
rect 31465 23745 31499 23773
rect 31527 23745 31561 23773
rect 31589 23745 31623 23773
rect 31651 23745 31699 23773
rect 31389 14959 31699 23745
rect 40264 23959 40424 23976
rect 40264 23931 40299 23959
rect 40327 23931 40361 23959
rect 40389 23931 40424 23959
rect 40264 23897 40424 23931
rect 40264 23869 40299 23897
rect 40327 23869 40361 23897
rect 40389 23869 40424 23897
rect 40264 23835 40424 23869
rect 40264 23807 40299 23835
rect 40327 23807 40361 23835
rect 40389 23807 40424 23835
rect 40264 23773 40424 23807
rect 40264 23745 40299 23773
rect 40327 23745 40361 23773
rect 40389 23745 40424 23773
rect 40264 23728 40424 23745
rect 55624 23959 55784 23976
rect 55624 23931 55659 23959
rect 55687 23931 55721 23959
rect 55749 23931 55784 23959
rect 55624 23897 55784 23931
rect 55624 23869 55659 23897
rect 55687 23869 55721 23897
rect 55749 23869 55784 23897
rect 55624 23835 55784 23869
rect 55624 23807 55659 23835
rect 55687 23807 55721 23835
rect 55749 23807 55784 23835
rect 55624 23773 55784 23807
rect 55624 23745 55659 23773
rect 55687 23745 55721 23773
rect 55749 23745 55784 23773
rect 55624 23728 55784 23745
rect 70984 23959 71144 23976
rect 70984 23931 71019 23959
rect 71047 23931 71081 23959
rect 71109 23931 71144 23959
rect 70984 23897 71144 23931
rect 70984 23869 71019 23897
rect 71047 23869 71081 23897
rect 71109 23869 71144 23897
rect 70984 23835 71144 23869
rect 70984 23807 71019 23835
rect 71047 23807 71081 23835
rect 71109 23807 71144 23835
rect 70984 23773 71144 23807
rect 70984 23745 71019 23773
rect 71047 23745 71081 23773
rect 71109 23745 71144 23773
rect 70984 23728 71144 23745
rect 86344 23959 86504 23976
rect 86344 23931 86379 23959
rect 86407 23931 86441 23959
rect 86469 23931 86504 23959
rect 86344 23897 86504 23931
rect 86344 23869 86379 23897
rect 86407 23869 86441 23897
rect 86469 23869 86504 23897
rect 86344 23835 86504 23869
rect 86344 23807 86379 23835
rect 86407 23807 86441 23835
rect 86469 23807 86504 23835
rect 86344 23773 86504 23807
rect 86344 23745 86379 23773
rect 86407 23745 86441 23773
rect 86469 23745 86504 23773
rect 86344 23728 86504 23745
rect 101704 23959 101864 23976
rect 101704 23931 101739 23959
rect 101767 23931 101801 23959
rect 101829 23931 101864 23959
rect 101704 23897 101864 23931
rect 101704 23869 101739 23897
rect 101767 23869 101801 23897
rect 101829 23869 101864 23897
rect 101704 23835 101864 23869
rect 101704 23807 101739 23835
rect 101767 23807 101801 23835
rect 101829 23807 101864 23835
rect 101704 23773 101864 23807
rect 101704 23745 101739 23773
rect 101767 23745 101801 23773
rect 101829 23745 101864 23773
rect 101704 23728 101864 23745
rect 117064 23959 117224 23976
rect 117064 23931 117099 23959
rect 117127 23931 117161 23959
rect 117189 23931 117224 23959
rect 117064 23897 117224 23931
rect 117064 23869 117099 23897
rect 117127 23869 117161 23897
rect 117189 23869 117224 23897
rect 117064 23835 117224 23869
rect 117064 23807 117099 23835
rect 117127 23807 117161 23835
rect 117189 23807 117224 23835
rect 117064 23773 117224 23807
rect 117064 23745 117099 23773
rect 117127 23745 117161 23773
rect 117189 23745 117224 23773
rect 117064 23728 117224 23745
rect 132424 23959 132584 23976
rect 132424 23931 132459 23959
rect 132487 23931 132521 23959
rect 132549 23931 132584 23959
rect 132424 23897 132584 23931
rect 132424 23869 132459 23897
rect 132487 23869 132521 23897
rect 132549 23869 132584 23897
rect 132424 23835 132584 23869
rect 132424 23807 132459 23835
rect 132487 23807 132521 23835
rect 132549 23807 132584 23835
rect 132424 23773 132584 23807
rect 132424 23745 132459 23773
rect 132487 23745 132521 23773
rect 132549 23745 132584 23773
rect 132424 23728 132584 23745
rect 147784 23959 147944 23976
rect 147784 23931 147819 23959
rect 147847 23931 147881 23959
rect 147909 23931 147944 23959
rect 147784 23897 147944 23931
rect 147784 23869 147819 23897
rect 147847 23869 147881 23897
rect 147909 23869 147944 23897
rect 147784 23835 147944 23869
rect 147784 23807 147819 23835
rect 147847 23807 147881 23835
rect 147909 23807 147944 23835
rect 147784 23773 147944 23807
rect 147784 23745 147819 23773
rect 147847 23745 147881 23773
rect 147909 23745 147944 23773
rect 147784 23728 147944 23745
rect 163144 23959 163304 23976
rect 163144 23931 163179 23959
rect 163207 23931 163241 23959
rect 163269 23931 163304 23959
rect 163144 23897 163304 23931
rect 163144 23869 163179 23897
rect 163207 23869 163241 23897
rect 163269 23869 163304 23897
rect 163144 23835 163304 23869
rect 163144 23807 163179 23835
rect 163207 23807 163241 23835
rect 163269 23807 163304 23835
rect 163144 23773 163304 23807
rect 163144 23745 163179 23773
rect 163207 23745 163241 23773
rect 163269 23745 163304 23773
rect 163144 23728 163304 23745
rect 178504 23959 178664 23976
rect 178504 23931 178539 23959
rect 178567 23931 178601 23959
rect 178629 23931 178664 23959
rect 178504 23897 178664 23931
rect 178504 23869 178539 23897
rect 178567 23869 178601 23897
rect 178629 23869 178664 23897
rect 178504 23835 178664 23869
rect 178504 23807 178539 23835
rect 178567 23807 178601 23835
rect 178629 23807 178664 23835
rect 178504 23773 178664 23807
rect 178504 23745 178539 23773
rect 178567 23745 178601 23773
rect 178629 23745 178664 23773
rect 178504 23728 178664 23745
rect 193864 23959 194024 23976
rect 193864 23931 193899 23959
rect 193927 23931 193961 23959
rect 193989 23931 194024 23959
rect 193864 23897 194024 23931
rect 193864 23869 193899 23897
rect 193927 23869 193961 23897
rect 193989 23869 194024 23897
rect 193864 23835 194024 23869
rect 193864 23807 193899 23835
rect 193927 23807 193961 23835
rect 193989 23807 194024 23835
rect 193864 23773 194024 23807
rect 193864 23745 193899 23773
rect 193927 23745 193961 23773
rect 193989 23745 194024 23773
rect 193864 23728 194024 23745
rect 209224 23959 209384 23976
rect 209224 23931 209259 23959
rect 209287 23931 209321 23959
rect 209349 23931 209384 23959
rect 209224 23897 209384 23931
rect 209224 23869 209259 23897
rect 209287 23869 209321 23897
rect 209349 23869 209384 23897
rect 209224 23835 209384 23869
rect 209224 23807 209259 23835
rect 209287 23807 209321 23835
rect 209349 23807 209384 23835
rect 209224 23773 209384 23807
rect 209224 23745 209259 23773
rect 209287 23745 209321 23773
rect 209349 23745 209384 23773
rect 209224 23728 209384 23745
rect 224584 23959 224744 23976
rect 224584 23931 224619 23959
rect 224647 23931 224681 23959
rect 224709 23931 224744 23959
rect 224584 23897 224744 23931
rect 224584 23869 224619 23897
rect 224647 23869 224681 23897
rect 224709 23869 224744 23897
rect 224584 23835 224744 23869
rect 224584 23807 224619 23835
rect 224647 23807 224681 23835
rect 224709 23807 224744 23835
rect 224584 23773 224744 23807
rect 224584 23745 224619 23773
rect 224647 23745 224681 23773
rect 224709 23745 224744 23773
rect 224584 23728 224744 23745
rect 239944 23959 240104 23976
rect 239944 23931 239979 23959
rect 240007 23931 240041 23959
rect 240069 23931 240104 23959
rect 239944 23897 240104 23931
rect 239944 23869 239979 23897
rect 240007 23869 240041 23897
rect 240069 23869 240104 23897
rect 239944 23835 240104 23869
rect 239944 23807 239979 23835
rect 240007 23807 240041 23835
rect 240069 23807 240104 23835
rect 239944 23773 240104 23807
rect 239944 23745 239979 23773
rect 240007 23745 240041 23773
rect 240069 23745 240104 23773
rect 239944 23728 240104 23745
rect 32584 20959 32744 20976
rect 32584 20931 32619 20959
rect 32647 20931 32681 20959
rect 32709 20931 32744 20959
rect 32584 20897 32744 20931
rect 32584 20869 32619 20897
rect 32647 20869 32681 20897
rect 32709 20869 32744 20897
rect 32584 20835 32744 20869
rect 32584 20807 32619 20835
rect 32647 20807 32681 20835
rect 32709 20807 32744 20835
rect 32584 20773 32744 20807
rect 32584 20745 32619 20773
rect 32647 20745 32681 20773
rect 32709 20745 32744 20773
rect 32584 20728 32744 20745
rect 47944 20959 48104 20976
rect 47944 20931 47979 20959
rect 48007 20931 48041 20959
rect 48069 20931 48104 20959
rect 47944 20897 48104 20931
rect 47944 20869 47979 20897
rect 48007 20869 48041 20897
rect 48069 20869 48104 20897
rect 47944 20835 48104 20869
rect 47944 20807 47979 20835
rect 48007 20807 48041 20835
rect 48069 20807 48104 20835
rect 47944 20773 48104 20807
rect 47944 20745 47979 20773
rect 48007 20745 48041 20773
rect 48069 20745 48104 20773
rect 47944 20728 48104 20745
rect 63304 20959 63464 20976
rect 63304 20931 63339 20959
rect 63367 20931 63401 20959
rect 63429 20931 63464 20959
rect 63304 20897 63464 20931
rect 63304 20869 63339 20897
rect 63367 20869 63401 20897
rect 63429 20869 63464 20897
rect 63304 20835 63464 20869
rect 63304 20807 63339 20835
rect 63367 20807 63401 20835
rect 63429 20807 63464 20835
rect 63304 20773 63464 20807
rect 63304 20745 63339 20773
rect 63367 20745 63401 20773
rect 63429 20745 63464 20773
rect 63304 20728 63464 20745
rect 78664 20959 78824 20976
rect 78664 20931 78699 20959
rect 78727 20931 78761 20959
rect 78789 20931 78824 20959
rect 78664 20897 78824 20931
rect 78664 20869 78699 20897
rect 78727 20869 78761 20897
rect 78789 20869 78824 20897
rect 78664 20835 78824 20869
rect 78664 20807 78699 20835
rect 78727 20807 78761 20835
rect 78789 20807 78824 20835
rect 78664 20773 78824 20807
rect 78664 20745 78699 20773
rect 78727 20745 78761 20773
rect 78789 20745 78824 20773
rect 78664 20728 78824 20745
rect 94024 20959 94184 20976
rect 94024 20931 94059 20959
rect 94087 20931 94121 20959
rect 94149 20931 94184 20959
rect 94024 20897 94184 20931
rect 94024 20869 94059 20897
rect 94087 20869 94121 20897
rect 94149 20869 94184 20897
rect 94024 20835 94184 20869
rect 94024 20807 94059 20835
rect 94087 20807 94121 20835
rect 94149 20807 94184 20835
rect 94024 20773 94184 20807
rect 94024 20745 94059 20773
rect 94087 20745 94121 20773
rect 94149 20745 94184 20773
rect 94024 20728 94184 20745
rect 109384 20959 109544 20976
rect 109384 20931 109419 20959
rect 109447 20931 109481 20959
rect 109509 20931 109544 20959
rect 109384 20897 109544 20931
rect 109384 20869 109419 20897
rect 109447 20869 109481 20897
rect 109509 20869 109544 20897
rect 109384 20835 109544 20869
rect 109384 20807 109419 20835
rect 109447 20807 109481 20835
rect 109509 20807 109544 20835
rect 109384 20773 109544 20807
rect 109384 20745 109419 20773
rect 109447 20745 109481 20773
rect 109509 20745 109544 20773
rect 109384 20728 109544 20745
rect 124744 20959 124904 20976
rect 124744 20931 124779 20959
rect 124807 20931 124841 20959
rect 124869 20931 124904 20959
rect 124744 20897 124904 20931
rect 124744 20869 124779 20897
rect 124807 20869 124841 20897
rect 124869 20869 124904 20897
rect 124744 20835 124904 20869
rect 124744 20807 124779 20835
rect 124807 20807 124841 20835
rect 124869 20807 124904 20835
rect 124744 20773 124904 20807
rect 124744 20745 124779 20773
rect 124807 20745 124841 20773
rect 124869 20745 124904 20773
rect 124744 20728 124904 20745
rect 140104 20959 140264 20976
rect 140104 20931 140139 20959
rect 140167 20931 140201 20959
rect 140229 20931 140264 20959
rect 140104 20897 140264 20931
rect 140104 20869 140139 20897
rect 140167 20869 140201 20897
rect 140229 20869 140264 20897
rect 140104 20835 140264 20869
rect 140104 20807 140139 20835
rect 140167 20807 140201 20835
rect 140229 20807 140264 20835
rect 140104 20773 140264 20807
rect 140104 20745 140139 20773
rect 140167 20745 140201 20773
rect 140229 20745 140264 20773
rect 140104 20728 140264 20745
rect 155464 20959 155624 20976
rect 155464 20931 155499 20959
rect 155527 20931 155561 20959
rect 155589 20931 155624 20959
rect 155464 20897 155624 20931
rect 155464 20869 155499 20897
rect 155527 20869 155561 20897
rect 155589 20869 155624 20897
rect 155464 20835 155624 20869
rect 155464 20807 155499 20835
rect 155527 20807 155561 20835
rect 155589 20807 155624 20835
rect 155464 20773 155624 20807
rect 155464 20745 155499 20773
rect 155527 20745 155561 20773
rect 155589 20745 155624 20773
rect 155464 20728 155624 20745
rect 170824 20959 170984 20976
rect 170824 20931 170859 20959
rect 170887 20931 170921 20959
rect 170949 20931 170984 20959
rect 170824 20897 170984 20931
rect 170824 20869 170859 20897
rect 170887 20869 170921 20897
rect 170949 20869 170984 20897
rect 170824 20835 170984 20869
rect 170824 20807 170859 20835
rect 170887 20807 170921 20835
rect 170949 20807 170984 20835
rect 170824 20773 170984 20807
rect 170824 20745 170859 20773
rect 170887 20745 170921 20773
rect 170949 20745 170984 20773
rect 170824 20728 170984 20745
rect 186184 20959 186344 20976
rect 186184 20931 186219 20959
rect 186247 20931 186281 20959
rect 186309 20931 186344 20959
rect 186184 20897 186344 20931
rect 186184 20869 186219 20897
rect 186247 20869 186281 20897
rect 186309 20869 186344 20897
rect 186184 20835 186344 20869
rect 186184 20807 186219 20835
rect 186247 20807 186281 20835
rect 186309 20807 186344 20835
rect 186184 20773 186344 20807
rect 186184 20745 186219 20773
rect 186247 20745 186281 20773
rect 186309 20745 186344 20773
rect 186184 20728 186344 20745
rect 201544 20959 201704 20976
rect 201544 20931 201579 20959
rect 201607 20931 201641 20959
rect 201669 20931 201704 20959
rect 201544 20897 201704 20931
rect 201544 20869 201579 20897
rect 201607 20869 201641 20897
rect 201669 20869 201704 20897
rect 201544 20835 201704 20869
rect 201544 20807 201579 20835
rect 201607 20807 201641 20835
rect 201669 20807 201704 20835
rect 201544 20773 201704 20807
rect 201544 20745 201579 20773
rect 201607 20745 201641 20773
rect 201669 20745 201704 20773
rect 201544 20728 201704 20745
rect 216904 20959 217064 20976
rect 216904 20931 216939 20959
rect 216967 20931 217001 20959
rect 217029 20931 217064 20959
rect 216904 20897 217064 20931
rect 216904 20869 216939 20897
rect 216967 20869 217001 20897
rect 217029 20869 217064 20897
rect 216904 20835 217064 20869
rect 216904 20807 216939 20835
rect 216967 20807 217001 20835
rect 217029 20807 217064 20835
rect 216904 20773 217064 20807
rect 216904 20745 216939 20773
rect 216967 20745 217001 20773
rect 217029 20745 217064 20773
rect 216904 20728 217064 20745
rect 232264 20959 232424 20976
rect 232264 20931 232299 20959
rect 232327 20931 232361 20959
rect 232389 20931 232424 20959
rect 232264 20897 232424 20931
rect 232264 20869 232299 20897
rect 232327 20869 232361 20897
rect 232389 20869 232424 20897
rect 232264 20835 232424 20869
rect 232264 20807 232299 20835
rect 232327 20807 232361 20835
rect 232389 20807 232424 20835
rect 232264 20773 232424 20807
rect 232264 20745 232299 20773
rect 232327 20745 232361 20773
rect 232389 20745 232424 20773
rect 232264 20728 232424 20745
rect 247624 20959 247784 20976
rect 247624 20931 247659 20959
rect 247687 20931 247721 20959
rect 247749 20931 247784 20959
rect 247624 20897 247784 20931
rect 247624 20869 247659 20897
rect 247687 20869 247721 20897
rect 247749 20869 247784 20897
rect 247624 20835 247784 20869
rect 247624 20807 247659 20835
rect 247687 20807 247721 20835
rect 247749 20807 247784 20835
rect 247624 20773 247784 20807
rect 247624 20745 247659 20773
rect 247687 20745 247721 20773
rect 247749 20745 247784 20773
rect 247624 20728 247784 20745
rect 254529 20959 254839 29745
rect 254529 20931 254577 20959
rect 254605 20931 254639 20959
rect 254667 20931 254701 20959
rect 254729 20931 254763 20959
rect 254791 20931 254839 20959
rect 254529 20897 254839 20931
rect 254529 20869 254577 20897
rect 254605 20869 254639 20897
rect 254667 20869 254701 20897
rect 254729 20869 254763 20897
rect 254791 20869 254839 20897
rect 254529 20835 254839 20869
rect 254529 20807 254577 20835
rect 254605 20807 254639 20835
rect 254667 20807 254701 20835
rect 254729 20807 254763 20835
rect 254791 20807 254839 20835
rect 254529 20773 254839 20807
rect 254529 20745 254577 20773
rect 254605 20745 254639 20773
rect 254667 20745 254701 20773
rect 254729 20745 254763 20773
rect 254791 20745 254839 20773
rect 31389 14931 31437 14959
rect 31465 14931 31499 14959
rect 31527 14931 31561 14959
rect 31589 14931 31623 14959
rect 31651 14931 31699 14959
rect 31389 14897 31699 14931
rect 31389 14869 31437 14897
rect 31465 14869 31499 14897
rect 31527 14869 31561 14897
rect 31589 14869 31623 14897
rect 31651 14869 31699 14897
rect 31389 14835 31699 14869
rect 31389 14807 31437 14835
rect 31465 14807 31499 14835
rect 31527 14807 31561 14835
rect 31589 14807 31623 14835
rect 31651 14807 31699 14835
rect 31389 14773 31699 14807
rect 31389 14745 31437 14773
rect 31465 14745 31499 14773
rect 31527 14745 31561 14773
rect 31589 14745 31623 14773
rect 31651 14745 31699 14773
rect 31389 5959 31699 14745
rect 247389 14959 247699 15510
rect 247389 14931 247437 14959
rect 247465 14931 247499 14959
rect 247527 14931 247561 14959
rect 247589 14931 247623 14959
rect 247651 14931 247699 14959
rect 247389 14897 247699 14931
rect 247389 14869 247437 14897
rect 247465 14869 247499 14897
rect 247527 14869 247561 14897
rect 247589 14869 247623 14897
rect 247651 14869 247699 14897
rect 247389 14835 247699 14869
rect 247389 14807 247437 14835
rect 247465 14807 247499 14835
rect 247527 14807 247561 14835
rect 247589 14807 247623 14835
rect 247651 14807 247699 14835
rect 247389 14773 247699 14807
rect 247389 14745 247437 14773
rect 247465 14745 247499 14773
rect 247527 14745 247561 14773
rect 247589 14745 247623 14773
rect 247651 14745 247699 14773
rect 31389 5931 31437 5959
rect 31465 5931 31499 5959
rect 31527 5931 31561 5959
rect 31589 5931 31623 5959
rect 31651 5931 31699 5959
rect 31389 5897 31699 5931
rect 31389 5869 31437 5897
rect 31465 5869 31499 5897
rect 31527 5869 31561 5897
rect 31589 5869 31623 5897
rect 31651 5869 31699 5897
rect 31389 5835 31699 5869
rect 31389 5807 31437 5835
rect 31465 5807 31499 5835
rect 31527 5807 31561 5835
rect 31589 5807 31623 5835
rect 31651 5807 31699 5835
rect 31389 5773 31699 5807
rect 31389 5745 31437 5773
rect 31465 5745 31499 5773
rect 31527 5745 31561 5773
rect 31589 5745 31623 5773
rect 31651 5745 31699 5773
rect 31389 424 31699 5745
rect 31389 396 31437 424
rect 31465 396 31499 424
rect 31527 396 31561 424
rect 31589 396 31623 424
rect 31651 396 31699 424
rect 31389 362 31699 396
rect 31389 334 31437 362
rect 31465 334 31499 362
rect 31527 334 31561 362
rect 31589 334 31623 362
rect 31651 334 31699 362
rect 31389 300 31699 334
rect 31389 272 31437 300
rect 31465 272 31499 300
rect 31527 272 31561 300
rect 31589 272 31623 300
rect 31651 272 31699 300
rect 31389 238 31699 272
rect 31389 210 31437 238
rect 31465 210 31499 238
rect 31527 210 31561 238
rect 31589 210 31623 238
rect 31651 210 31699 238
rect 31389 162 31699 210
rect 38529 11959 38839 14541
rect 38529 11931 38577 11959
rect 38605 11931 38639 11959
rect 38667 11931 38701 11959
rect 38729 11931 38763 11959
rect 38791 11931 38839 11959
rect 38529 11897 38839 11931
rect 38529 11869 38577 11897
rect 38605 11869 38639 11897
rect 38667 11869 38701 11897
rect 38729 11869 38763 11897
rect 38791 11869 38839 11897
rect 38529 11835 38839 11869
rect 38529 11807 38577 11835
rect 38605 11807 38639 11835
rect 38667 11807 38701 11835
rect 38729 11807 38763 11835
rect 38791 11807 38839 11835
rect 38529 11773 38839 11807
rect 38529 11745 38577 11773
rect 38605 11745 38639 11773
rect 38667 11745 38701 11773
rect 38729 11745 38763 11773
rect 38791 11745 38839 11773
rect 38529 2959 38839 11745
rect 38529 2931 38577 2959
rect 38605 2931 38639 2959
rect 38667 2931 38701 2959
rect 38729 2931 38763 2959
rect 38791 2931 38839 2959
rect 38529 2897 38839 2931
rect 38529 2869 38577 2897
rect 38605 2869 38639 2897
rect 38667 2869 38701 2897
rect 38729 2869 38763 2897
rect 38791 2869 38839 2897
rect 38529 2835 38839 2869
rect 38529 2807 38577 2835
rect 38605 2807 38639 2835
rect 38667 2807 38701 2835
rect 38729 2807 38763 2835
rect 38791 2807 38839 2835
rect 38529 2773 38839 2807
rect 38529 2745 38577 2773
rect 38605 2745 38639 2773
rect 38667 2745 38701 2773
rect 38729 2745 38763 2773
rect 38791 2745 38839 2773
rect 38529 904 38839 2745
rect 38529 876 38577 904
rect 38605 876 38639 904
rect 38667 876 38701 904
rect 38729 876 38763 904
rect 38791 876 38839 904
rect 38529 842 38839 876
rect 38529 814 38577 842
rect 38605 814 38639 842
rect 38667 814 38701 842
rect 38729 814 38763 842
rect 38791 814 38839 842
rect 38529 780 38839 814
rect 38529 752 38577 780
rect 38605 752 38639 780
rect 38667 752 38701 780
rect 38729 752 38763 780
rect 38791 752 38839 780
rect 38529 718 38839 752
rect 38529 690 38577 718
rect 38605 690 38639 718
rect 38667 690 38701 718
rect 38729 690 38763 718
rect 38791 690 38839 718
rect 38529 162 38839 690
rect 40389 5959 40699 14541
rect 40389 5931 40437 5959
rect 40465 5931 40499 5959
rect 40527 5931 40561 5959
rect 40589 5931 40623 5959
rect 40651 5931 40699 5959
rect 40389 5897 40699 5931
rect 40389 5869 40437 5897
rect 40465 5869 40499 5897
rect 40527 5869 40561 5897
rect 40589 5869 40623 5897
rect 40651 5869 40699 5897
rect 40389 5835 40699 5869
rect 40389 5807 40437 5835
rect 40465 5807 40499 5835
rect 40527 5807 40561 5835
rect 40589 5807 40623 5835
rect 40651 5807 40699 5835
rect 40389 5773 40699 5807
rect 40389 5745 40437 5773
rect 40465 5745 40499 5773
rect 40527 5745 40561 5773
rect 40589 5745 40623 5773
rect 40651 5745 40699 5773
rect 40389 424 40699 5745
rect 40389 396 40437 424
rect 40465 396 40499 424
rect 40527 396 40561 424
rect 40589 396 40623 424
rect 40651 396 40699 424
rect 40389 362 40699 396
rect 40389 334 40437 362
rect 40465 334 40499 362
rect 40527 334 40561 362
rect 40589 334 40623 362
rect 40651 334 40699 362
rect 40389 300 40699 334
rect 40389 272 40437 300
rect 40465 272 40499 300
rect 40527 272 40561 300
rect 40589 272 40623 300
rect 40651 272 40699 300
rect 40389 238 40699 272
rect 40389 210 40437 238
rect 40465 210 40499 238
rect 40527 210 40561 238
rect 40589 210 40623 238
rect 40651 210 40699 238
rect 40389 162 40699 210
rect 47529 11959 47839 14541
rect 47529 11931 47577 11959
rect 47605 11931 47639 11959
rect 47667 11931 47701 11959
rect 47729 11931 47763 11959
rect 47791 11931 47839 11959
rect 47529 11897 47839 11931
rect 47529 11869 47577 11897
rect 47605 11869 47639 11897
rect 47667 11869 47701 11897
rect 47729 11869 47763 11897
rect 47791 11869 47839 11897
rect 47529 11835 47839 11869
rect 47529 11807 47577 11835
rect 47605 11807 47639 11835
rect 47667 11807 47701 11835
rect 47729 11807 47763 11835
rect 47791 11807 47839 11835
rect 47529 11773 47839 11807
rect 47529 11745 47577 11773
rect 47605 11745 47639 11773
rect 47667 11745 47701 11773
rect 47729 11745 47763 11773
rect 47791 11745 47839 11773
rect 47529 2959 47839 11745
rect 47529 2931 47577 2959
rect 47605 2931 47639 2959
rect 47667 2931 47701 2959
rect 47729 2931 47763 2959
rect 47791 2931 47839 2959
rect 47529 2897 47839 2931
rect 47529 2869 47577 2897
rect 47605 2869 47639 2897
rect 47667 2869 47701 2897
rect 47729 2869 47763 2897
rect 47791 2869 47839 2897
rect 47529 2835 47839 2869
rect 47529 2807 47577 2835
rect 47605 2807 47639 2835
rect 47667 2807 47701 2835
rect 47729 2807 47763 2835
rect 47791 2807 47839 2835
rect 47529 2773 47839 2807
rect 47529 2745 47577 2773
rect 47605 2745 47639 2773
rect 47667 2745 47701 2773
rect 47729 2745 47763 2773
rect 47791 2745 47839 2773
rect 47529 904 47839 2745
rect 47529 876 47577 904
rect 47605 876 47639 904
rect 47667 876 47701 904
rect 47729 876 47763 904
rect 47791 876 47839 904
rect 47529 842 47839 876
rect 47529 814 47577 842
rect 47605 814 47639 842
rect 47667 814 47701 842
rect 47729 814 47763 842
rect 47791 814 47839 842
rect 47529 780 47839 814
rect 47529 752 47577 780
rect 47605 752 47639 780
rect 47667 752 47701 780
rect 47729 752 47763 780
rect 47791 752 47839 780
rect 47529 718 47839 752
rect 47529 690 47577 718
rect 47605 690 47639 718
rect 47667 690 47701 718
rect 47729 690 47763 718
rect 47791 690 47839 718
rect 47529 162 47839 690
rect 49389 5959 49699 14541
rect 49389 5931 49437 5959
rect 49465 5931 49499 5959
rect 49527 5931 49561 5959
rect 49589 5931 49623 5959
rect 49651 5931 49699 5959
rect 49389 5897 49699 5931
rect 49389 5869 49437 5897
rect 49465 5869 49499 5897
rect 49527 5869 49561 5897
rect 49589 5869 49623 5897
rect 49651 5869 49699 5897
rect 49389 5835 49699 5869
rect 49389 5807 49437 5835
rect 49465 5807 49499 5835
rect 49527 5807 49561 5835
rect 49589 5807 49623 5835
rect 49651 5807 49699 5835
rect 49389 5773 49699 5807
rect 49389 5745 49437 5773
rect 49465 5745 49499 5773
rect 49527 5745 49561 5773
rect 49589 5745 49623 5773
rect 49651 5745 49699 5773
rect 49389 424 49699 5745
rect 49389 396 49437 424
rect 49465 396 49499 424
rect 49527 396 49561 424
rect 49589 396 49623 424
rect 49651 396 49699 424
rect 49389 362 49699 396
rect 49389 334 49437 362
rect 49465 334 49499 362
rect 49527 334 49561 362
rect 49589 334 49623 362
rect 49651 334 49699 362
rect 49389 300 49699 334
rect 49389 272 49437 300
rect 49465 272 49499 300
rect 49527 272 49561 300
rect 49589 272 49623 300
rect 49651 272 49699 300
rect 49389 238 49699 272
rect 49389 210 49437 238
rect 49465 210 49499 238
rect 49527 210 49561 238
rect 49589 210 49623 238
rect 49651 210 49699 238
rect 49389 162 49699 210
rect 56529 11959 56839 14541
rect 56529 11931 56577 11959
rect 56605 11931 56639 11959
rect 56667 11931 56701 11959
rect 56729 11931 56763 11959
rect 56791 11931 56839 11959
rect 56529 11897 56839 11931
rect 56529 11869 56577 11897
rect 56605 11869 56639 11897
rect 56667 11869 56701 11897
rect 56729 11869 56763 11897
rect 56791 11869 56839 11897
rect 56529 11835 56839 11869
rect 56529 11807 56577 11835
rect 56605 11807 56639 11835
rect 56667 11807 56701 11835
rect 56729 11807 56763 11835
rect 56791 11807 56839 11835
rect 56529 11773 56839 11807
rect 56529 11745 56577 11773
rect 56605 11745 56639 11773
rect 56667 11745 56701 11773
rect 56729 11745 56763 11773
rect 56791 11745 56839 11773
rect 56529 2959 56839 11745
rect 56529 2931 56577 2959
rect 56605 2931 56639 2959
rect 56667 2931 56701 2959
rect 56729 2931 56763 2959
rect 56791 2931 56839 2959
rect 56529 2897 56839 2931
rect 56529 2869 56577 2897
rect 56605 2869 56639 2897
rect 56667 2869 56701 2897
rect 56729 2869 56763 2897
rect 56791 2869 56839 2897
rect 56529 2835 56839 2869
rect 56529 2807 56577 2835
rect 56605 2807 56639 2835
rect 56667 2807 56701 2835
rect 56729 2807 56763 2835
rect 56791 2807 56839 2835
rect 56529 2773 56839 2807
rect 56529 2745 56577 2773
rect 56605 2745 56639 2773
rect 56667 2745 56701 2773
rect 56729 2745 56763 2773
rect 56791 2745 56839 2773
rect 56529 904 56839 2745
rect 56529 876 56577 904
rect 56605 876 56639 904
rect 56667 876 56701 904
rect 56729 876 56763 904
rect 56791 876 56839 904
rect 56529 842 56839 876
rect 56529 814 56577 842
rect 56605 814 56639 842
rect 56667 814 56701 842
rect 56729 814 56763 842
rect 56791 814 56839 842
rect 56529 780 56839 814
rect 56529 752 56577 780
rect 56605 752 56639 780
rect 56667 752 56701 780
rect 56729 752 56763 780
rect 56791 752 56839 780
rect 56529 718 56839 752
rect 56529 690 56577 718
rect 56605 690 56639 718
rect 56667 690 56701 718
rect 56729 690 56763 718
rect 56791 690 56839 718
rect 56529 162 56839 690
rect 58389 5959 58699 14541
rect 58389 5931 58437 5959
rect 58465 5931 58499 5959
rect 58527 5931 58561 5959
rect 58589 5931 58623 5959
rect 58651 5931 58699 5959
rect 58389 5897 58699 5931
rect 58389 5869 58437 5897
rect 58465 5869 58499 5897
rect 58527 5869 58561 5897
rect 58589 5869 58623 5897
rect 58651 5869 58699 5897
rect 58389 5835 58699 5869
rect 58389 5807 58437 5835
rect 58465 5807 58499 5835
rect 58527 5807 58561 5835
rect 58589 5807 58623 5835
rect 58651 5807 58699 5835
rect 58389 5773 58699 5807
rect 58389 5745 58437 5773
rect 58465 5745 58499 5773
rect 58527 5745 58561 5773
rect 58589 5745 58623 5773
rect 58651 5745 58699 5773
rect 58389 424 58699 5745
rect 58389 396 58437 424
rect 58465 396 58499 424
rect 58527 396 58561 424
rect 58589 396 58623 424
rect 58651 396 58699 424
rect 58389 362 58699 396
rect 58389 334 58437 362
rect 58465 334 58499 362
rect 58527 334 58561 362
rect 58589 334 58623 362
rect 58651 334 58699 362
rect 58389 300 58699 334
rect 58389 272 58437 300
rect 58465 272 58499 300
rect 58527 272 58561 300
rect 58589 272 58623 300
rect 58651 272 58699 300
rect 58389 238 58699 272
rect 58389 210 58437 238
rect 58465 210 58499 238
rect 58527 210 58561 238
rect 58589 210 58623 238
rect 58651 210 58699 238
rect 58389 162 58699 210
rect 65529 11959 65839 14541
rect 65529 11931 65577 11959
rect 65605 11931 65639 11959
rect 65667 11931 65701 11959
rect 65729 11931 65763 11959
rect 65791 11931 65839 11959
rect 65529 11897 65839 11931
rect 65529 11869 65577 11897
rect 65605 11869 65639 11897
rect 65667 11869 65701 11897
rect 65729 11869 65763 11897
rect 65791 11869 65839 11897
rect 65529 11835 65839 11869
rect 65529 11807 65577 11835
rect 65605 11807 65639 11835
rect 65667 11807 65701 11835
rect 65729 11807 65763 11835
rect 65791 11807 65839 11835
rect 65529 11773 65839 11807
rect 65529 11745 65577 11773
rect 65605 11745 65639 11773
rect 65667 11745 65701 11773
rect 65729 11745 65763 11773
rect 65791 11745 65839 11773
rect 65529 2959 65839 11745
rect 65529 2931 65577 2959
rect 65605 2931 65639 2959
rect 65667 2931 65701 2959
rect 65729 2931 65763 2959
rect 65791 2931 65839 2959
rect 65529 2897 65839 2931
rect 65529 2869 65577 2897
rect 65605 2869 65639 2897
rect 65667 2869 65701 2897
rect 65729 2869 65763 2897
rect 65791 2869 65839 2897
rect 65529 2835 65839 2869
rect 65529 2807 65577 2835
rect 65605 2807 65639 2835
rect 65667 2807 65701 2835
rect 65729 2807 65763 2835
rect 65791 2807 65839 2835
rect 65529 2773 65839 2807
rect 65529 2745 65577 2773
rect 65605 2745 65639 2773
rect 65667 2745 65701 2773
rect 65729 2745 65763 2773
rect 65791 2745 65839 2773
rect 65529 904 65839 2745
rect 65529 876 65577 904
rect 65605 876 65639 904
rect 65667 876 65701 904
rect 65729 876 65763 904
rect 65791 876 65839 904
rect 65529 842 65839 876
rect 65529 814 65577 842
rect 65605 814 65639 842
rect 65667 814 65701 842
rect 65729 814 65763 842
rect 65791 814 65839 842
rect 65529 780 65839 814
rect 65529 752 65577 780
rect 65605 752 65639 780
rect 65667 752 65701 780
rect 65729 752 65763 780
rect 65791 752 65839 780
rect 65529 718 65839 752
rect 65529 690 65577 718
rect 65605 690 65639 718
rect 65667 690 65701 718
rect 65729 690 65763 718
rect 65791 690 65839 718
rect 65529 162 65839 690
rect 67389 5959 67699 14541
rect 67389 5931 67437 5959
rect 67465 5931 67499 5959
rect 67527 5931 67561 5959
rect 67589 5931 67623 5959
rect 67651 5931 67699 5959
rect 67389 5897 67699 5931
rect 67389 5869 67437 5897
rect 67465 5869 67499 5897
rect 67527 5869 67561 5897
rect 67589 5869 67623 5897
rect 67651 5869 67699 5897
rect 67389 5835 67699 5869
rect 67389 5807 67437 5835
rect 67465 5807 67499 5835
rect 67527 5807 67561 5835
rect 67589 5807 67623 5835
rect 67651 5807 67699 5835
rect 67389 5773 67699 5807
rect 67389 5745 67437 5773
rect 67465 5745 67499 5773
rect 67527 5745 67561 5773
rect 67589 5745 67623 5773
rect 67651 5745 67699 5773
rect 67389 424 67699 5745
rect 67389 396 67437 424
rect 67465 396 67499 424
rect 67527 396 67561 424
rect 67589 396 67623 424
rect 67651 396 67699 424
rect 67389 362 67699 396
rect 67389 334 67437 362
rect 67465 334 67499 362
rect 67527 334 67561 362
rect 67589 334 67623 362
rect 67651 334 67699 362
rect 67389 300 67699 334
rect 67389 272 67437 300
rect 67465 272 67499 300
rect 67527 272 67561 300
rect 67589 272 67623 300
rect 67651 272 67699 300
rect 67389 238 67699 272
rect 67389 210 67437 238
rect 67465 210 67499 238
rect 67527 210 67561 238
rect 67589 210 67623 238
rect 67651 210 67699 238
rect 67389 162 67699 210
rect 74529 11959 74839 14541
rect 74529 11931 74577 11959
rect 74605 11931 74639 11959
rect 74667 11931 74701 11959
rect 74729 11931 74763 11959
rect 74791 11931 74839 11959
rect 74529 11897 74839 11931
rect 74529 11869 74577 11897
rect 74605 11869 74639 11897
rect 74667 11869 74701 11897
rect 74729 11869 74763 11897
rect 74791 11869 74839 11897
rect 74529 11835 74839 11869
rect 74529 11807 74577 11835
rect 74605 11807 74639 11835
rect 74667 11807 74701 11835
rect 74729 11807 74763 11835
rect 74791 11807 74839 11835
rect 74529 11773 74839 11807
rect 74529 11745 74577 11773
rect 74605 11745 74639 11773
rect 74667 11745 74701 11773
rect 74729 11745 74763 11773
rect 74791 11745 74839 11773
rect 74529 2959 74839 11745
rect 74529 2931 74577 2959
rect 74605 2931 74639 2959
rect 74667 2931 74701 2959
rect 74729 2931 74763 2959
rect 74791 2931 74839 2959
rect 74529 2897 74839 2931
rect 74529 2869 74577 2897
rect 74605 2869 74639 2897
rect 74667 2869 74701 2897
rect 74729 2869 74763 2897
rect 74791 2869 74839 2897
rect 74529 2835 74839 2869
rect 74529 2807 74577 2835
rect 74605 2807 74639 2835
rect 74667 2807 74701 2835
rect 74729 2807 74763 2835
rect 74791 2807 74839 2835
rect 74529 2773 74839 2807
rect 74529 2745 74577 2773
rect 74605 2745 74639 2773
rect 74667 2745 74701 2773
rect 74729 2745 74763 2773
rect 74791 2745 74839 2773
rect 74529 904 74839 2745
rect 74529 876 74577 904
rect 74605 876 74639 904
rect 74667 876 74701 904
rect 74729 876 74763 904
rect 74791 876 74839 904
rect 74529 842 74839 876
rect 74529 814 74577 842
rect 74605 814 74639 842
rect 74667 814 74701 842
rect 74729 814 74763 842
rect 74791 814 74839 842
rect 74529 780 74839 814
rect 74529 752 74577 780
rect 74605 752 74639 780
rect 74667 752 74701 780
rect 74729 752 74763 780
rect 74791 752 74839 780
rect 74529 718 74839 752
rect 74529 690 74577 718
rect 74605 690 74639 718
rect 74667 690 74701 718
rect 74729 690 74763 718
rect 74791 690 74839 718
rect 74529 162 74839 690
rect 76389 5959 76699 14541
rect 76389 5931 76437 5959
rect 76465 5931 76499 5959
rect 76527 5931 76561 5959
rect 76589 5931 76623 5959
rect 76651 5931 76699 5959
rect 76389 5897 76699 5931
rect 76389 5869 76437 5897
rect 76465 5869 76499 5897
rect 76527 5869 76561 5897
rect 76589 5869 76623 5897
rect 76651 5869 76699 5897
rect 76389 5835 76699 5869
rect 76389 5807 76437 5835
rect 76465 5807 76499 5835
rect 76527 5807 76561 5835
rect 76589 5807 76623 5835
rect 76651 5807 76699 5835
rect 76389 5773 76699 5807
rect 76389 5745 76437 5773
rect 76465 5745 76499 5773
rect 76527 5745 76561 5773
rect 76589 5745 76623 5773
rect 76651 5745 76699 5773
rect 76389 424 76699 5745
rect 76389 396 76437 424
rect 76465 396 76499 424
rect 76527 396 76561 424
rect 76589 396 76623 424
rect 76651 396 76699 424
rect 76389 362 76699 396
rect 76389 334 76437 362
rect 76465 334 76499 362
rect 76527 334 76561 362
rect 76589 334 76623 362
rect 76651 334 76699 362
rect 76389 300 76699 334
rect 76389 272 76437 300
rect 76465 272 76499 300
rect 76527 272 76561 300
rect 76589 272 76623 300
rect 76651 272 76699 300
rect 76389 238 76699 272
rect 76389 210 76437 238
rect 76465 210 76499 238
rect 76527 210 76561 238
rect 76589 210 76623 238
rect 76651 210 76699 238
rect 76389 162 76699 210
rect 83529 11959 83839 14541
rect 83529 11931 83577 11959
rect 83605 11931 83639 11959
rect 83667 11931 83701 11959
rect 83729 11931 83763 11959
rect 83791 11931 83839 11959
rect 83529 11897 83839 11931
rect 83529 11869 83577 11897
rect 83605 11869 83639 11897
rect 83667 11869 83701 11897
rect 83729 11869 83763 11897
rect 83791 11869 83839 11897
rect 83529 11835 83839 11869
rect 83529 11807 83577 11835
rect 83605 11807 83639 11835
rect 83667 11807 83701 11835
rect 83729 11807 83763 11835
rect 83791 11807 83839 11835
rect 83529 11773 83839 11807
rect 83529 11745 83577 11773
rect 83605 11745 83639 11773
rect 83667 11745 83701 11773
rect 83729 11745 83763 11773
rect 83791 11745 83839 11773
rect 83529 2959 83839 11745
rect 83529 2931 83577 2959
rect 83605 2931 83639 2959
rect 83667 2931 83701 2959
rect 83729 2931 83763 2959
rect 83791 2931 83839 2959
rect 83529 2897 83839 2931
rect 83529 2869 83577 2897
rect 83605 2869 83639 2897
rect 83667 2869 83701 2897
rect 83729 2869 83763 2897
rect 83791 2869 83839 2897
rect 83529 2835 83839 2869
rect 83529 2807 83577 2835
rect 83605 2807 83639 2835
rect 83667 2807 83701 2835
rect 83729 2807 83763 2835
rect 83791 2807 83839 2835
rect 83529 2773 83839 2807
rect 83529 2745 83577 2773
rect 83605 2745 83639 2773
rect 83667 2745 83701 2773
rect 83729 2745 83763 2773
rect 83791 2745 83839 2773
rect 83529 904 83839 2745
rect 83529 876 83577 904
rect 83605 876 83639 904
rect 83667 876 83701 904
rect 83729 876 83763 904
rect 83791 876 83839 904
rect 83529 842 83839 876
rect 83529 814 83577 842
rect 83605 814 83639 842
rect 83667 814 83701 842
rect 83729 814 83763 842
rect 83791 814 83839 842
rect 83529 780 83839 814
rect 83529 752 83577 780
rect 83605 752 83639 780
rect 83667 752 83701 780
rect 83729 752 83763 780
rect 83791 752 83839 780
rect 83529 718 83839 752
rect 83529 690 83577 718
rect 83605 690 83639 718
rect 83667 690 83701 718
rect 83729 690 83763 718
rect 83791 690 83839 718
rect 83529 162 83839 690
rect 85389 5959 85699 14541
rect 85389 5931 85437 5959
rect 85465 5931 85499 5959
rect 85527 5931 85561 5959
rect 85589 5931 85623 5959
rect 85651 5931 85699 5959
rect 85389 5897 85699 5931
rect 85389 5869 85437 5897
rect 85465 5869 85499 5897
rect 85527 5869 85561 5897
rect 85589 5869 85623 5897
rect 85651 5869 85699 5897
rect 85389 5835 85699 5869
rect 85389 5807 85437 5835
rect 85465 5807 85499 5835
rect 85527 5807 85561 5835
rect 85589 5807 85623 5835
rect 85651 5807 85699 5835
rect 85389 5773 85699 5807
rect 85389 5745 85437 5773
rect 85465 5745 85499 5773
rect 85527 5745 85561 5773
rect 85589 5745 85623 5773
rect 85651 5745 85699 5773
rect 85389 424 85699 5745
rect 85389 396 85437 424
rect 85465 396 85499 424
rect 85527 396 85561 424
rect 85589 396 85623 424
rect 85651 396 85699 424
rect 85389 362 85699 396
rect 85389 334 85437 362
rect 85465 334 85499 362
rect 85527 334 85561 362
rect 85589 334 85623 362
rect 85651 334 85699 362
rect 85389 300 85699 334
rect 85389 272 85437 300
rect 85465 272 85499 300
rect 85527 272 85561 300
rect 85589 272 85623 300
rect 85651 272 85699 300
rect 85389 238 85699 272
rect 85389 210 85437 238
rect 85465 210 85499 238
rect 85527 210 85561 238
rect 85589 210 85623 238
rect 85651 210 85699 238
rect 85389 162 85699 210
rect 92529 11959 92839 14541
rect 92529 11931 92577 11959
rect 92605 11931 92639 11959
rect 92667 11931 92701 11959
rect 92729 11931 92763 11959
rect 92791 11931 92839 11959
rect 92529 11897 92839 11931
rect 92529 11869 92577 11897
rect 92605 11869 92639 11897
rect 92667 11869 92701 11897
rect 92729 11869 92763 11897
rect 92791 11869 92839 11897
rect 92529 11835 92839 11869
rect 92529 11807 92577 11835
rect 92605 11807 92639 11835
rect 92667 11807 92701 11835
rect 92729 11807 92763 11835
rect 92791 11807 92839 11835
rect 92529 11773 92839 11807
rect 92529 11745 92577 11773
rect 92605 11745 92639 11773
rect 92667 11745 92701 11773
rect 92729 11745 92763 11773
rect 92791 11745 92839 11773
rect 92529 2959 92839 11745
rect 92529 2931 92577 2959
rect 92605 2931 92639 2959
rect 92667 2931 92701 2959
rect 92729 2931 92763 2959
rect 92791 2931 92839 2959
rect 92529 2897 92839 2931
rect 92529 2869 92577 2897
rect 92605 2869 92639 2897
rect 92667 2869 92701 2897
rect 92729 2869 92763 2897
rect 92791 2869 92839 2897
rect 92529 2835 92839 2869
rect 92529 2807 92577 2835
rect 92605 2807 92639 2835
rect 92667 2807 92701 2835
rect 92729 2807 92763 2835
rect 92791 2807 92839 2835
rect 92529 2773 92839 2807
rect 92529 2745 92577 2773
rect 92605 2745 92639 2773
rect 92667 2745 92701 2773
rect 92729 2745 92763 2773
rect 92791 2745 92839 2773
rect 92529 904 92839 2745
rect 92529 876 92577 904
rect 92605 876 92639 904
rect 92667 876 92701 904
rect 92729 876 92763 904
rect 92791 876 92839 904
rect 92529 842 92839 876
rect 92529 814 92577 842
rect 92605 814 92639 842
rect 92667 814 92701 842
rect 92729 814 92763 842
rect 92791 814 92839 842
rect 92529 780 92839 814
rect 92529 752 92577 780
rect 92605 752 92639 780
rect 92667 752 92701 780
rect 92729 752 92763 780
rect 92791 752 92839 780
rect 92529 718 92839 752
rect 92529 690 92577 718
rect 92605 690 92639 718
rect 92667 690 92701 718
rect 92729 690 92763 718
rect 92791 690 92839 718
rect 92529 162 92839 690
rect 94389 5959 94699 14541
rect 94389 5931 94437 5959
rect 94465 5931 94499 5959
rect 94527 5931 94561 5959
rect 94589 5931 94623 5959
rect 94651 5931 94699 5959
rect 94389 5897 94699 5931
rect 94389 5869 94437 5897
rect 94465 5869 94499 5897
rect 94527 5869 94561 5897
rect 94589 5869 94623 5897
rect 94651 5869 94699 5897
rect 94389 5835 94699 5869
rect 94389 5807 94437 5835
rect 94465 5807 94499 5835
rect 94527 5807 94561 5835
rect 94589 5807 94623 5835
rect 94651 5807 94699 5835
rect 94389 5773 94699 5807
rect 94389 5745 94437 5773
rect 94465 5745 94499 5773
rect 94527 5745 94561 5773
rect 94589 5745 94623 5773
rect 94651 5745 94699 5773
rect 94389 424 94699 5745
rect 94389 396 94437 424
rect 94465 396 94499 424
rect 94527 396 94561 424
rect 94589 396 94623 424
rect 94651 396 94699 424
rect 94389 362 94699 396
rect 94389 334 94437 362
rect 94465 334 94499 362
rect 94527 334 94561 362
rect 94589 334 94623 362
rect 94651 334 94699 362
rect 94389 300 94699 334
rect 94389 272 94437 300
rect 94465 272 94499 300
rect 94527 272 94561 300
rect 94589 272 94623 300
rect 94651 272 94699 300
rect 94389 238 94699 272
rect 94389 210 94437 238
rect 94465 210 94499 238
rect 94527 210 94561 238
rect 94589 210 94623 238
rect 94651 210 94699 238
rect 94389 162 94699 210
rect 101529 11959 101839 14541
rect 101529 11931 101577 11959
rect 101605 11931 101639 11959
rect 101667 11931 101701 11959
rect 101729 11931 101763 11959
rect 101791 11931 101839 11959
rect 101529 11897 101839 11931
rect 101529 11869 101577 11897
rect 101605 11869 101639 11897
rect 101667 11869 101701 11897
rect 101729 11869 101763 11897
rect 101791 11869 101839 11897
rect 101529 11835 101839 11869
rect 101529 11807 101577 11835
rect 101605 11807 101639 11835
rect 101667 11807 101701 11835
rect 101729 11807 101763 11835
rect 101791 11807 101839 11835
rect 101529 11773 101839 11807
rect 101529 11745 101577 11773
rect 101605 11745 101639 11773
rect 101667 11745 101701 11773
rect 101729 11745 101763 11773
rect 101791 11745 101839 11773
rect 101529 2959 101839 11745
rect 101529 2931 101577 2959
rect 101605 2931 101639 2959
rect 101667 2931 101701 2959
rect 101729 2931 101763 2959
rect 101791 2931 101839 2959
rect 101529 2897 101839 2931
rect 101529 2869 101577 2897
rect 101605 2869 101639 2897
rect 101667 2869 101701 2897
rect 101729 2869 101763 2897
rect 101791 2869 101839 2897
rect 101529 2835 101839 2869
rect 101529 2807 101577 2835
rect 101605 2807 101639 2835
rect 101667 2807 101701 2835
rect 101729 2807 101763 2835
rect 101791 2807 101839 2835
rect 101529 2773 101839 2807
rect 101529 2745 101577 2773
rect 101605 2745 101639 2773
rect 101667 2745 101701 2773
rect 101729 2745 101763 2773
rect 101791 2745 101839 2773
rect 101529 904 101839 2745
rect 101529 876 101577 904
rect 101605 876 101639 904
rect 101667 876 101701 904
rect 101729 876 101763 904
rect 101791 876 101839 904
rect 101529 842 101839 876
rect 101529 814 101577 842
rect 101605 814 101639 842
rect 101667 814 101701 842
rect 101729 814 101763 842
rect 101791 814 101839 842
rect 101529 780 101839 814
rect 101529 752 101577 780
rect 101605 752 101639 780
rect 101667 752 101701 780
rect 101729 752 101763 780
rect 101791 752 101839 780
rect 101529 718 101839 752
rect 101529 690 101577 718
rect 101605 690 101639 718
rect 101667 690 101701 718
rect 101729 690 101763 718
rect 101791 690 101839 718
rect 101529 162 101839 690
rect 103389 5959 103699 14541
rect 103389 5931 103437 5959
rect 103465 5931 103499 5959
rect 103527 5931 103561 5959
rect 103589 5931 103623 5959
rect 103651 5931 103699 5959
rect 103389 5897 103699 5931
rect 103389 5869 103437 5897
rect 103465 5869 103499 5897
rect 103527 5869 103561 5897
rect 103589 5869 103623 5897
rect 103651 5869 103699 5897
rect 103389 5835 103699 5869
rect 103389 5807 103437 5835
rect 103465 5807 103499 5835
rect 103527 5807 103561 5835
rect 103589 5807 103623 5835
rect 103651 5807 103699 5835
rect 103389 5773 103699 5807
rect 103389 5745 103437 5773
rect 103465 5745 103499 5773
rect 103527 5745 103561 5773
rect 103589 5745 103623 5773
rect 103651 5745 103699 5773
rect 103389 424 103699 5745
rect 103389 396 103437 424
rect 103465 396 103499 424
rect 103527 396 103561 424
rect 103589 396 103623 424
rect 103651 396 103699 424
rect 103389 362 103699 396
rect 103389 334 103437 362
rect 103465 334 103499 362
rect 103527 334 103561 362
rect 103589 334 103623 362
rect 103651 334 103699 362
rect 103389 300 103699 334
rect 103389 272 103437 300
rect 103465 272 103499 300
rect 103527 272 103561 300
rect 103589 272 103623 300
rect 103651 272 103699 300
rect 103389 238 103699 272
rect 103389 210 103437 238
rect 103465 210 103499 238
rect 103527 210 103561 238
rect 103589 210 103623 238
rect 103651 210 103699 238
rect 103389 162 103699 210
rect 110529 11959 110839 14541
rect 110529 11931 110577 11959
rect 110605 11931 110639 11959
rect 110667 11931 110701 11959
rect 110729 11931 110763 11959
rect 110791 11931 110839 11959
rect 110529 11897 110839 11931
rect 110529 11869 110577 11897
rect 110605 11869 110639 11897
rect 110667 11869 110701 11897
rect 110729 11869 110763 11897
rect 110791 11869 110839 11897
rect 110529 11835 110839 11869
rect 110529 11807 110577 11835
rect 110605 11807 110639 11835
rect 110667 11807 110701 11835
rect 110729 11807 110763 11835
rect 110791 11807 110839 11835
rect 110529 11773 110839 11807
rect 110529 11745 110577 11773
rect 110605 11745 110639 11773
rect 110667 11745 110701 11773
rect 110729 11745 110763 11773
rect 110791 11745 110839 11773
rect 110529 2959 110839 11745
rect 110529 2931 110577 2959
rect 110605 2931 110639 2959
rect 110667 2931 110701 2959
rect 110729 2931 110763 2959
rect 110791 2931 110839 2959
rect 110529 2897 110839 2931
rect 110529 2869 110577 2897
rect 110605 2869 110639 2897
rect 110667 2869 110701 2897
rect 110729 2869 110763 2897
rect 110791 2869 110839 2897
rect 110529 2835 110839 2869
rect 110529 2807 110577 2835
rect 110605 2807 110639 2835
rect 110667 2807 110701 2835
rect 110729 2807 110763 2835
rect 110791 2807 110839 2835
rect 110529 2773 110839 2807
rect 110529 2745 110577 2773
rect 110605 2745 110639 2773
rect 110667 2745 110701 2773
rect 110729 2745 110763 2773
rect 110791 2745 110839 2773
rect 110529 904 110839 2745
rect 110529 876 110577 904
rect 110605 876 110639 904
rect 110667 876 110701 904
rect 110729 876 110763 904
rect 110791 876 110839 904
rect 110529 842 110839 876
rect 110529 814 110577 842
rect 110605 814 110639 842
rect 110667 814 110701 842
rect 110729 814 110763 842
rect 110791 814 110839 842
rect 110529 780 110839 814
rect 110529 752 110577 780
rect 110605 752 110639 780
rect 110667 752 110701 780
rect 110729 752 110763 780
rect 110791 752 110839 780
rect 110529 718 110839 752
rect 110529 690 110577 718
rect 110605 690 110639 718
rect 110667 690 110701 718
rect 110729 690 110763 718
rect 110791 690 110839 718
rect 110529 162 110839 690
rect 112389 5959 112699 14541
rect 112389 5931 112437 5959
rect 112465 5931 112499 5959
rect 112527 5931 112561 5959
rect 112589 5931 112623 5959
rect 112651 5931 112699 5959
rect 112389 5897 112699 5931
rect 112389 5869 112437 5897
rect 112465 5869 112499 5897
rect 112527 5869 112561 5897
rect 112589 5869 112623 5897
rect 112651 5869 112699 5897
rect 112389 5835 112699 5869
rect 112389 5807 112437 5835
rect 112465 5807 112499 5835
rect 112527 5807 112561 5835
rect 112589 5807 112623 5835
rect 112651 5807 112699 5835
rect 112389 5773 112699 5807
rect 112389 5745 112437 5773
rect 112465 5745 112499 5773
rect 112527 5745 112561 5773
rect 112589 5745 112623 5773
rect 112651 5745 112699 5773
rect 112389 424 112699 5745
rect 112389 396 112437 424
rect 112465 396 112499 424
rect 112527 396 112561 424
rect 112589 396 112623 424
rect 112651 396 112699 424
rect 112389 362 112699 396
rect 112389 334 112437 362
rect 112465 334 112499 362
rect 112527 334 112561 362
rect 112589 334 112623 362
rect 112651 334 112699 362
rect 112389 300 112699 334
rect 112389 272 112437 300
rect 112465 272 112499 300
rect 112527 272 112561 300
rect 112589 272 112623 300
rect 112651 272 112699 300
rect 112389 238 112699 272
rect 112389 210 112437 238
rect 112465 210 112499 238
rect 112527 210 112561 238
rect 112589 210 112623 238
rect 112651 210 112699 238
rect 112389 162 112699 210
rect 119529 11959 119839 14541
rect 119529 11931 119577 11959
rect 119605 11931 119639 11959
rect 119667 11931 119701 11959
rect 119729 11931 119763 11959
rect 119791 11931 119839 11959
rect 119529 11897 119839 11931
rect 119529 11869 119577 11897
rect 119605 11869 119639 11897
rect 119667 11869 119701 11897
rect 119729 11869 119763 11897
rect 119791 11869 119839 11897
rect 119529 11835 119839 11869
rect 119529 11807 119577 11835
rect 119605 11807 119639 11835
rect 119667 11807 119701 11835
rect 119729 11807 119763 11835
rect 119791 11807 119839 11835
rect 119529 11773 119839 11807
rect 119529 11745 119577 11773
rect 119605 11745 119639 11773
rect 119667 11745 119701 11773
rect 119729 11745 119763 11773
rect 119791 11745 119839 11773
rect 119529 2959 119839 11745
rect 119529 2931 119577 2959
rect 119605 2931 119639 2959
rect 119667 2931 119701 2959
rect 119729 2931 119763 2959
rect 119791 2931 119839 2959
rect 119529 2897 119839 2931
rect 119529 2869 119577 2897
rect 119605 2869 119639 2897
rect 119667 2869 119701 2897
rect 119729 2869 119763 2897
rect 119791 2869 119839 2897
rect 119529 2835 119839 2869
rect 119529 2807 119577 2835
rect 119605 2807 119639 2835
rect 119667 2807 119701 2835
rect 119729 2807 119763 2835
rect 119791 2807 119839 2835
rect 119529 2773 119839 2807
rect 119529 2745 119577 2773
rect 119605 2745 119639 2773
rect 119667 2745 119701 2773
rect 119729 2745 119763 2773
rect 119791 2745 119839 2773
rect 119529 904 119839 2745
rect 119529 876 119577 904
rect 119605 876 119639 904
rect 119667 876 119701 904
rect 119729 876 119763 904
rect 119791 876 119839 904
rect 119529 842 119839 876
rect 119529 814 119577 842
rect 119605 814 119639 842
rect 119667 814 119701 842
rect 119729 814 119763 842
rect 119791 814 119839 842
rect 119529 780 119839 814
rect 119529 752 119577 780
rect 119605 752 119639 780
rect 119667 752 119701 780
rect 119729 752 119763 780
rect 119791 752 119839 780
rect 119529 718 119839 752
rect 119529 690 119577 718
rect 119605 690 119639 718
rect 119667 690 119701 718
rect 119729 690 119763 718
rect 119791 690 119839 718
rect 119529 162 119839 690
rect 121389 5959 121699 14541
rect 121389 5931 121437 5959
rect 121465 5931 121499 5959
rect 121527 5931 121561 5959
rect 121589 5931 121623 5959
rect 121651 5931 121699 5959
rect 121389 5897 121699 5931
rect 121389 5869 121437 5897
rect 121465 5869 121499 5897
rect 121527 5869 121561 5897
rect 121589 5869 121623 5897
rect 121651 5869 121699 5897
rect 121389 5835 121699 5869
rect 121389 5807 121437 5835
rect 121465 5807 121499 5835
rect 121527 5807 121561 5835
rect 121589 5807 121623 5835
rect 121651 5807 121699 5835
rect 121389 5773 121699 5807
rect 121389 5745 121437 5773
rect 121465 5745 121499 5773
rect 121527 5745 121561 5773
rect 121589 5745 121623 5773
rect 121651 5745 121699 5773
rect 121389 424 121699 5745
rect 121389 396 121437 424
rect 121465 396 121499 424
rect 121527 396 121561 424
rect 121589 396 121623 424
rect 121651 396 121699 424
rect 121389 362 121699 396
rect 121389 334 121437 362
rect 121465 334 121499 362
rect 121527 334 121561 362
rect 121589 334 121623 362
rect 121651 334 121699 362
rect 121389 300 121699 334
rect 121389 272 121437 300
rect 121465 272 121499 300
rect 121527 272 121561 300
rect 121589 272 121623 300
rect 121651 272 121699 300
rect 121389 238 121699 272
rect 121389 210 121437 238
rect 121465 210 121499 238
rect 121527 210 121561 238
rect 121589 210 121623 238
rect 121651 210 121699 238
rect 121389 162 121699 210
rect 128529 11959 128839 14541
rect 128529 11931 128577 11959
rect 128605 11931 128639 11959
rect 128667 11931 128701 11959
rect 128729 11931 128763 11959
rect 128791 11931 128839 11959
rect 128529 11897 128839 11931
rect 128529 11869 128577 11897
rect 128605 11869 128639 11897
rect 128667 11869 128701 11897
rect 128729 11869 128763 11897
rect 128791 11869 128839 11897
rect 128529 11835 128839 11869
rect 128529 11807 128577 11835
rect 128605 11807 128639 11835
rect 128667 11807 128701 11835
rect 128729 11807 128763 11835
rect 128791 11807 128839 11835
rect 128529 11773 128839 11807
rect 128529 11745 128577 11773
rect 128605 11745 128639 11773
rect 128667 11745 128701 11773
rect 128729 11745 128763 11773
rect 128791 11745 128839 11773
rect 128529 2959 128839 11745
rect 128529 2931 128577 2959
rect 128605 2931 128639 2959
rect 128667 2931 128701 2959
rect 128729 2931 128763 2959
rect 128791 2931 128839 2959
rect 128529 2897 128839 2931
rect 128529 2869 128577 2897
rect 128605 2869 128639 2897
rect 128667 2869 128701 2897
rect 128729 2869 128763 2897
rect 128791 2869 128839 2897
rect 128529 2835 128839 2869
rect 128529 2807 128577 2835
rect 128605 2807 128639 2835
rect 128667 2807 128701 2835
rect 128729 2807 128763 2835
rect 128791 2807 128839 2835
rect 128529 2773 128839 2807
rect 128529 2745 128577 2773
rect 128605 2745 128639 2773
rect 128667 2745 128701 2773
rect 128729 2745 128763 2773
rect 128791 2745 128839 2773
rect 128529 904 128839 2745
rect 128529 876 128577 904
rect 128605 876 128639 904
rect 128667 876 128701 904
rect 128729 876 128763 904
rect 128791 876 128839 904
rect 128529 842 128839 876
rect 128529 814 128577 842
rect 128605 814 128639 842
rect 128667 814 128701 842
rect 128729 814 128763 842
rect 128791 814 128839 842
rect 128529 780 128839 814
rect 128529 752 128577 780
rect 128605 752 128639 780
rect 128667 752 128701 780
rect 128729 752 128763 780
rect 128791 752 128839 780
rect 128529 718 128839 752
rect 128529 690 128577 718
rect 128605 690 128639 718
rect 128667 690 128701 718
rect 128729 690 128763 718
rect 128791 690 128839 718
rect 128529 162 128839 690
rect 130389 5959 130699 14541
rect 130389 5931 130437 5959
rect 130465 5931 130499 5959
rect 130527 5931 130561 5959
rect 130589 5931 130623 5959
rect 130651 5931 130699 5959
rect 130389 5897 130699 5931
rect 130389 5869 130437 5897
rect 130465 5869 130499 5897
rect 130527 5869 130561 5897
rect 130589 5869 130623 5897
rect 130651 5869 130699 5897
rect 130389 5835 130699 5869
rect 130389 5807 130437 5835
rect 130465 5807 130499 5835
rect 130527 5807 130561 5835
rect 130589 5807 130623 5835
rect 130651 5807 130699 5835
rect 130389 5773 130699 5807
rect 130389 5745 130437 5773
rect 130465 5745 130499 5773
rect 130527 5745 130561 5773
rect 130589 5745 130623 5773
rect 130651 5745 130699 5773
rect 130389 424 130699 5745
rect 130389 396 130437 424
rect 130465 396 130499 424
rect 130527 396 130561 424
rect 130589 396 130623 424
rect 130651 396 130699 424
rect 130389 362 130699 396
rect 130389 334 130437 362
rect 130465 334 130499 362
rect 130527 334 130561 362
rect 130589 334 130623 362
rect 130651 334 130699 362
rect 130389 300 130699 334
rect 130389 272 130437 300
rect 130465 272 130499 300
rect 130527 272 130561 300
rect 130589 272 130623 300
rect 130651 272 130699 300
rect 130389 238 130699 272
rect 130389 210 130437 238
rect 130465 210 130499 238
rect 130527 210 130561 238
rect 130589 210 130623 238
rect 130651 210 130699 238
rect 130389 162 130699 210
rect 137529 11959 137839 14541
rect 137529 11931 137577 11959
rect 137605 11931 137639 11959
rect 137667 11931 137701 11959
rect 137729 11931 137763 11959
rect 137791 11931 137839 11959
rect 137529 11897 137839 11931
rect 137529 11869 137577 11897
rect 137605 11869 137639 11897
rect 137667 11869 137701 11897
rect 137729 11869 137763 11897
rect 137791 11869 137839 11897
rect 137529 11835 137839 11869
rect 137529 11807 137577 11835
rect 137605 11807 137639 11835
rect 137667 11807 137701 11835
rect 137729 11807 137763 11835
rect 137791 11807 137839 11835
rect 137529 11773 137839 11807
rect 137529 11745 137577 11773
rect 137605 11745 137639 11773
rect 137667 11745 137701 11773
rect 137729 11745 137763 11773
rect 137791 11745 137839 11773
rect 137529 2959 137839 11745
rect 137529 2931 137577 2959
rect 137605 2931 137639 2959
rect 137667 2931 137701 2959
rect 137729 2931 137763 2959
rect 137791 2931 137839 2959
rect 137529 2897 137839 2931
rect 137529 2869 137577 2897
rect 137605 2869 137639 2897
rect 137667 2869 137701 2897
rect 137729 2869 137763 2897
rect 137791 2869 137839 2897
rect 137529 2835 137839 2869
rect 137529 2807 137577 2835
rect 137605 2807 137639 2835
rect 137667 2807 137701 2835
rect 137729 2807 137763 2835
rect 137791 2807 137839 2835
rect 137529 2773 137839 2807
rect 137529 2745 137577 2773
rect 137605 2745 137639 2773
rect 137667 2745 137701 2773
rect 137729 2745 137763 2773
rect 137791 2745 137839 2773
rect 137529 904 137839 2745
rect 137529 876 137577 904
rect 137605 876 137639 904
rect 137667 876 137701 904
rect 137729 876 137763 904
rect 137791 876 137839 904
rect 137529 842 137839 876
rect 137529 814 137577 842
rect 137605 814 137639 842
rect 137667 814 137701 842
rect 137729 814 137763 842
rect 137791 814 137839 842
rect 137529 780 137839 814
rect 137529 752 137577 780
rect 137605 752 137639 780
rect 137667 752 137701 780
rect 137729 752 137763 780
rect 137791 752 137839 780
rect 137529 718 137839 752
rect 137529 690 137577 718
rect 137605 690 137639 718
rect 137667 690 137701 718
rect 137729 690 137763 718
rect 137791 690 137839 718
rect 137529 162 137839 690
rect 139389 5959 139699 14541
rect 139389 5931 139437 5959
rect 139465 5931 139499 5959
rect 139527 5931 139561 5959
rect 139589 5931 139623 5959
rect 139651 5931 139699 5959
rect 139389 5897 139699 5931
rect 139389 5869 139437 5897
rect 139465 5869 139499 5897
rect 139527 5869 139561 5897
rect 139589 5869 139623 5897
rect 139651 5869 139699 5897
rect 139389 5835 139699 5869
rect 139389 5807 139437 5835
rect 139465 5807 139499 5835
rect 139527 5807 139561 5835
rect 139589 5807 139623 5835
rect 139651 5807 139699 5835
rect 139389 5773 139699 5807
rect 139389 5745 139437 5773
rect 139465 5745 139499 5773
rect 139527 5745 139561 5773
rect 139589 5745 139623 5773
rect 139651 5745 139699 5773
rect 139389 424 139699 5745
rect 139389 396 139437 424
rect 139465 396 139499 424
rect 139527 396 139561 424
rect 139589 396 139623 424
rect 139651 396 139699 424
rect 139389 362 139699 396
rect 139389 334 139437 362
rect 139465 334 139499 362
rect 139527 334 139561 362
rect 139589 334 139623 362
rect 139651 334 139699 362
rect 139389 300 139699 334
rect 139389 272 139437 300
rect 139465 272 139499 300
rect 139527 272 139561 300
rect 139589 272 139623 300
rect 139651 272 139699 300
rect 139389 238 139699 272
rect 139389 210 139437 238
rect 139465 210 139499 238
rect 139527 210 139561 238
rect 139589 210 139623 238
rect 139651 210 139699 238
rect 139389 162 139699 210
rect 146529 11959 146839 14541
rect 146529 11931 146577 11959
rect 146605 11931 146639 11959
rect 146667 11931 146701 11959
rect 146729 11931 146763 11959
rect 146791 11931 146839 11959
rect 146529 11897 146839 11931
rect 146529 11869 146577 11897
rect 146605 11869 146639 11897
rect 146667 11869 146701 11897
rect 146729 11869 146763 11897
rect 146791 11869 146839 11897
rect 146529 11835 146839 11869
rect 146529 11807 146577 11835
rect 146605 11807 146639 11835
rect 146667 11807 146701 11835
rect 146729 11807 146763 11835
rect 146791 11807 146839 11835
rect 146529 11773 146839 11807
rect 146529 11745 146577 11773
rect 146605 11745 146639 11773
rect 146667 11745 146701 11773
rect 146729 11745 146763 11773
rect 146791 11745 146839 11773
rect 146529 2959 146839 11745
rect 146529 2931 146577 2959
rect 146605 2931 146639 2959
rect 146667 2931 146701 2959
rect 146729 2931 146763 2959
rect 146791 2931 146839 2959
rect 146529 2897 146839 2931
rect 146529 2869 146577 2897
rect 146605 2869 146639 2897
rect 146667 2869 146701 2897
rect 146729 2869 146763 2897
rect 146791 2869 146839 2897
rect 146529 2835 146839 2869
rect 146529 2807 146577 2835
rect 146605 2807 146639 2835
rect 146667 2807 146701 2835
rect 146729 2807 146763 2835
rect 146791 2807 146839 2835
rect 146529 2773 146839 2807
rect 146529 2745 146577 2773
rect 146605 2745 146639 2773
rect 146667 2745 146701 2773
rect 146729 2745 146763 2773
rect 146791 2745 146839 2773
rect 146529 904 146839 2745
rect 146529 876 146577 904
rect 146605 876 146639 904
rect 146667 876 146701 904
rect 146729 876 146763 904
rect 146791 876 146839 904
rect 146529 842 146839 876
rect 146529 814 146577 842
rect 146605 814 146639 842
rect 146667 814 146701 842
rect 146729 814 146763 842
rect 146791 814 146839 842
rect 146529 780 146839 814
rect 146529 752 146577 780
rect 146605 752 146639 780
rect 146667 752 146701 780
rect 146729 752 146763 780
rect 146791 752 146839 780
rect 146529 718 146839 752
rect 146529 690 146577 718
rect 146605 690 146639 718
rect 146667 690 146701 718
rect 146729 690 146763 718
rect 146791 690 146839 718
rect 146529 162 146839 690
rect 148389 5959 148699 14541
rect 148389 5931 148437 5959
rect 148465 5931 148499 5959
rect 148527 5931 148561 5959
rect 148589 5931 148623 5959
rect 148651 5931 148699 5959
rect 148389 5897 148699 5931
rect 148389 5869 148437 5897
rect 148465 5869 148499 5897
rect 148527 5869 148561 5897
rect 148589 5869 148623 5897
rect 148651 5869 148699 5897
rect 148389 5835 148699 5869
rect 148389 5807 148437 5835
rect 148465 5807 148499 5835
rect 148527 5807 148561 5835
rect 148589 5807 148623 5835
rect 148651 5807 148699 5835
rect 148389 5773 148699 5807
rect 148389 5745 148437 5773
rect 148465 5745 148499 5773
rect 148527 5745 148561 5773
rect 148589 5745 148623 5773
rect 148651 5745 148699 5773
rect 148389 424 148699 5745
rect 148389 396 148437 424
rect 148465 396 148499 424
rect 148527 396 148561 424
rect 148589 396 148623 424
rect 148651 396 148699 424
rect 148389 362 148699 396
rect 148389 334 148437 362
rect 148465 334 148499 362
rect 148527 334 148561 362
rect 148589 334 148623 362
rect 148651 334 148699 362
rect 148389 300 148699 334
rect 148389 272 148437 300
rect 148465 272 148499 300
rect 148527 272 148561 300
rect 148589 272 148623 300
rect 148651 272 148699 300
rect 148389 238 148699 272
rect 148389 210 148437 238
rect 148465 210 148499 238
rect 148527 210 148561 238
rect 148589 210 148623 238
rect 148651 210 148699 238
rect 148389 162 148699 210
rect 155529 11959 155839 14541
rect 155529 11931 155577 11959
rect 155605 11931 155639 11959
rect 155667 11931 155701 11959
rect 155729 11931 155763 11959
rect 155791 11931 155839 11959
rect 155529 11897 155839 11931
rect 155529 11869 155577 11897
rect 155605 11869 155639 11897
rect 155667 11869 155701 11897
rect 155729 11869 155763 11897
rect 155791 11869 155839 11897
rect 155529 11835 155839 11869
rect 155529 11807 155577 11835
rect 155605 11807 155639 11835
rect 155667 11807 155701 11835
rect 155729 11807 155763 11835
rect 155791 11807 155839 11835
rect 155529 11773 155839 11807
rect 155529 11745 155577 11773
rect 155605 11745 155639 11773
rect 155667 11745 155701 11773
rect 155729 11745 155763 11773
rect 155791 11745 155839 11773
rect 155529 2959 155839 11745
rect 155529 2931 155577 2959
rect 155605 2931 155639 2959
rect 155667 2931 155701 2959
rect 155729 2931 155763 2959
rect 155791 2931 155839 2959
rect 155529 2897 155839 2931
rect 155529 2869 155577 2897
rect 155605 2869 155639 2897
rect 155667 2869 155701 2897
rect 155729 2869 155763 2897
rect 155791 2869 155839 2897
rect 155529 2835 155839 2869
rect 155529 2807 155577 2835
rect 155605 2807 155639 2835
rect 155667 2807 155701 2835
rect 155729 2807 155763 2835
rect 155791 2807 155839 2835
rect 155529 2773 155839 2807
rect 155529 2745 155577 2773
rect 155605 2745 155639 2773
rect 155667 2745 155701 2773
rect 155729 2745 155763 2773
rect 155791 2745 155839 2773
rect 155529 904 155839 2745
rect 155529 876 155577 904
rect 155605 876 155639 904
rect 155667 876 155701 904
rect 155729 876 155763 904
rect 155791 876 155839 904
rect 155529 842 155839 876
rect 155529 814 155577 842
rect 155605 814 155639 842
rect 155667 814 155701 842
rect 155729 814 155763 842
rect 155791 814 155839 842
rect 155529 780 155839 814
rect 155529 752 155577 780
rect 155605 752 155639 780
rect 155667 752 155701 780
rect 155729 752 155763 780
rect 155791 752 155839 780
rect 155529 718 155839 752
rect 155529 690 155577 718
rect 155605 690 155639 718
rect 155667 690 155701 718
rect 155729 690 155763 718
rect 155791 690 155839 718
rect 155529 162 155839 690
rect 157389 5959 157699 14541
rect 157389 5931 157437 5959
rect 157465 5931 157499 5959
rect 157527 5931 157561 5959
rect 157589 5931 157623 5959
rect 157651 5931 157699 5959
rect 157389 5897 157699 5931
rect 157389 5869 157437 5897
rect 157465 5869 157499 5897
rect 157527 5869 157561 5897
rect 157589 5869 157623 5897
rect 157651 5869 157699 5897
rect 157389 5835 157699 5869
rect 157389 5807 157437 5835
rect 157465 5807 157499 5835
rect 157527 5807 157561 5835
rect 157589 5807 157623 5835
rect 157651 5807 157699 5835
rect 157389 5773 157699 5807
rect 157389 5745 157437 5773
rect 157465 5745 157499 5773
rect 157527 5745 157561 5773
rect 157589 5745 157623 5773
rect 157651 5745 157699 5773
rect 157389 424 157699 5745
rect 157389 396 157437 424
rect 157465 396 157499 424
rect 157527 396 157561 424
rect 157589 396 157623 424
rect 157651 396 157699 424
rect 157389 362 157699 396
rect 157389 334 157437 362
rect 157465 334 157499 362
rect 157527 334 157561 362
rect 157589 334 157623 362
rect 157651 334 157699 362
rect 157389 300 157699 334
rect 157389 272 157437 300
rect 157465 272 157499 300
rect 157527 272 157561 300
rect 157589 272 157623 300
rect 157651 272 157699 300
rect 157389 238 157699 272
rect 157389 210 157437 238
rect 157465 210 157499 238
rect 157527 210 157561 238
rect 157589 210 157623 238
rect 157651 210 157699 238
rect 157389 162 157699 210
rect 164529 11959 164839 14541
rect 164529 11931 164577 11959
rect 164605 11931 164639 11959
rect 164667 11931 164701 11959
rect 164729 11931 164763 11959
rect 164791 11931 164839 11959
rect 164529 11897 164839 11931
rect 164529 11869 164577 11897
rect 164605 11869 164639 11897
rect 164667 11869 164701 11897
rect 164729 11869 164763 11897
rect 164791 11869 164839 11897
rect 164529 11835 164839 11869
rect 164529 11807 164577 11835
rect 164605 11807 164639 11835
rect 164667 11807 164701 11835
rect 164729 11807 164763 11835
rect 164791 11807 164839 11835
rect 164529 11773 164839 11807
rect 164529 11745 164577 11773
rect 164605 11745 164639 11773
rect 164667 11745 164701 11773
rect 164729 11745 164763 11773
rect 164791 11745 164839 11773
rect 164529 2959 164839 11745
rect 164529 2931 164577 2959
rect 164605 2931 164639 2959
rect 164667 2931 164701 2959
rect 164729 2931 164763 2959
rect 164791 2931 164839 2959
rect 164529 2897 164839 2931
rect 164529 2869 164577 2897
rect 164605 2869 164639 2897
rect 164667 2869 164701 2897
rect 164729 2869 164763 2897
rect 164791 2869 164839 2897
rect 164529 2835 164839 2869
rect 164529 2807 164577 2835
rect 164605 2807 164639 2835
rect 164667 2807 164701 2835
rect 164729 2807 164763 2835
rect 164791 2807 164839 2835
rect 164529 2773 164839 2807
rect 164529 2745 164577 2773
rect 164605 2745 164639 2773
rect 164667 2745 164701 2773
rect 164729 2745 164763 2773
rect 164791 2745 164839 2773
rect 164529 904 164839 2745
rect 164529 876 164577 904
rect 164605 876 164639 904
rect 164667 876 164701 904
rect 164729 876 164763 904
rect 164791 876 164839 904
rect 164529 842 164839 876
rect 164529 814 164577 842
rect 164605 814 164639 842
rect 164667 814 164701 842
rect 164729 814 164763 842
rect 164791 814 164839 842
rect 164529 780 164839 814
rect 164529 752 164577 780
rect 164605 752 164639 780
rect 164667 752 164701 780
rect 164729 752 164763 780
rect 164791 752 164839 780
rect 164529 718 164839 752
rect 164529 690 164577 718
rect 164605 690 164639 718
rect 164667 690 164701 718
rect 164729 690 164763 718
rect 164791 690 164839 718
rect 164529 162 164839 690
rect 166389 5959 166699 14541
rect 166389 5931 166437 5959
rect 166465 5931 166499 5959
rect 166527 5931 166561 5959
rect 166589 5931 166623 5959
rect 166651 5931 166699 5959
rect 166389 5897 166699 5931
rect 166389 5869 166437 5897
rect 166465 5869 166499 5897
rect 166527 5869 166561 5897
rect 166589 5869 166623 5897
rect 166651 5869 166699 5897
rect 166389 5835 166699 5869
rect 166389 5807 166437 5835
rect 166465 5807 166499 5835
rect 166527 5807 166561 5835
rect 166589 5807 166623 5835
rect 166651 5807 166699 5835
rect 166389 5773 166699 5807
rect 166389 5745 166437 5773
rect 166465 5745 166499 5773
rect 166527 5745 166561 5773
rect 166589 5745 166623 5773
rect 166651 5745 166699 5773
rect 166389 424 166699 5745
rect 166389 396 166437 424
rect 166465 396 166499 424
rect 166527 396 166561 424
rect 166589 396 166623 424
rect 166651 396 166699 424
rect 166389 362 166699 396
rect 166389 334 166437 362
rect 166465 334 166499 362
rect 166527 334 166561 362
rect 166589 334 166623 362
rect 166651 334 166699 362
rect 166389 300 166699 334
rect 166389 272 166437 300
rect 166465 272 166499 300
rect 166527 272 166561 300
rect 166589 272 166623 300
rect 166651 272 166699 300
rect 166389 238 166699 272
rect 166389 210 166437 238
rect 166465 210 166499 238
rect 166527 210 166561 238
rect 166589 210 166623 238
rect 166651 210 166699 238
rect 166389 162 166699 210
rect 173529 11959 173839 14541
rect 173529 11931 173577 11959
rect 173605 11931 173639 11959
rect 173667 11931 173701 11959
rect 173729 11931 173763 11959
rect 173791 11931 173839 11959
rect 173529 11897 173839 11931
rect 173529 11869 173577 11897
rect 173605 11869 173639 11897
rect 173667 11869 173701 11897
rect 173729 11869 173763 11897
rect 173791 11869 173839 11897
rect 173529 11835 173839 11869
rect 173529 11807 173577 11835
rect 173605 11807 173639 11835
rect 173667 11807 173701 11835
rect 173729 11807 173763 11835
rect 173791 11807 173839 11835
rect 173529 11773 173839 11807
rect 173529 11745 173577 11773
rect 173605 11745 173639 11773
rect 173667 11745 173701 11773
rect 173729 11745 173763 11773
rect 173791 11745 173839 11773
rect 173529 2959 173839 11745
rect 173529 2931 173577 2959
rect 173605 2931 173639 2959
rect 173667 2931 173701 2959
rect 173729 2931 173763 2959
rect 173791 2931 173839 2959
rect 173529 2897 173839 2931
rect 173529 2869 173577 2897
rect 173605 2869 173639 2897
rect 173667 2869 173701 2897
rect 173729 2869 173763 2897
rect 173791 2869 173839 2897
rect 173529 2835 173839 2869
rect 173529 2807 173577 2835
rect 173605 2807 173639 2835
rect 173667 2807 173701 2835
rect 173729 2807 173763 2835
rect 173791 2807 173839 2835
rect 173529 2773 173839 2807
rect 173529 2745 173577 2773
rect 173605 2745 173639 2773
rect 173667 2745 173701 2773
rect 173729 2745 173763 2773
rect 173791 2745 173839 2773
rect 173529 904 173839 2745
rect 173529 876 173577 904
rect 173605 876 173639 904
rect 173667 876 173701 904
rect 173729 876 173763 904
rect 173791 876 173839 904
rect 173529 842 173839 876
rect 173529 814 173577 842
rect 173605 814 173639 842
rect 173667 814 173701 842
rect 173729 814 173763 842
rect 173791 814 173839 842
rect 173529 780 173839 814
rect 173529 752 173577 780
rect 173605 752 173639 780
rect 173667 752 173701 780
rect 173729 752 173763 780
rect 173791 752 173839 780
rect 173529 718 173839 752
rect 173529 690 173577 718
rect 173605 690 173639 718
rect 173667 690 173701 718
rect 173729 690 173763 718
rect 173791 690 173839 718
rect 173529 162 173839 690
rect 175389 5959 175699 14541
rect 175389 5931 175437 5959
rect 175465 5931 175499 5959
rect 175527 5931 175561 5959
rect 175589 5931 175623 5959
rect 175651 5931 175699 5959
rect 175389 5897 175699 5931
rect 175389 5869 175437 5897
rect 175465 5869 175499 5897
rect 175527 5869 175561 5897
rect 175589 5869 175623 5897
rect 175651 5869 175699 5897
rect 175389 5835 175699 5869
rect 175389 5807 175437 5835
rect 175465 5807 175499 5835
rect 175527 5807 175561 5835
rect 175589 5807 175623 5835
rect 175651 5807 175699 5835
rect 175389 5773 175699 5807
rect 175389 5745 175437 5773
rect 175465 5745 175499 5773
rect 175527 5745 175561 5773
rect 175589 5745 175623 5773
rect 175651 5745 175699 5773
rect 175389 424 175699 5745
rect 175389 396 175437 424
rect 175465 396 175499 424
rect 175527 396 175561 424
rect 175589 396 175623 424
rect 175651 396 175699 424
rect 175389 362 175699 396
rect 175389 334 175437 362
rect 175465 334 175499 362
rect 175527 334 175561 362
rect 175589 334 175623 362
rect 175651 334 175699 362
rect 175389 300 175699 334
rect 175389 272 175437 300
rect 175465 272 175499 300
rect 175527 272 175561 300
rect 175589 272 175623 300
rect 175651 272 175699 300
rect 175389 238 175699 272
rect 175389 210 175437 238
rect 175465 210 175499 238
rect 175527 210 175561 238
rect 175589 210 175623 238
rect 175651 210 175699 238
rect 175389 162 175699 210
rect 182529 11959 182839 14541
rect 182529 11931 182577 11959
rect 182605 11931 182639 11959
rect 182667 11931 182701 11959
rect 182729 11931 182763 11959
rect 182791 11931 182839 11959
rect 182529 11897 182839 11931
rect 182529 11869 182577 11897
rect 182605 11869 182639 11897
rect 182667 11869 182701 11897
rect 182729 11869 182763 11897
rect 182791 11869 182839 11897
rect 182529 11835 182839 11869
rect 182529 11807 182577 11835
rect 182605 11807 182639 11835
rect 182667 11807 182701 11835
rect 182729 11807 182763 11835
rect 182791 11807 182839 11835
rect 182529 11773 182839 11807
rect 182529 11745 182577 11773
rect 182605 11745 182639 11773
rect 182667 11745 182701 11773
rect 182729 11745 182763 11773
rect 182791 11745 182839 11773
rect 182529 2959 182839 11745
rect 182529 2931 182577 2959
rect 182605 2931 182639 2959
rect 182667 2931 182701 2959
rect 182729 2931 182763 2959
rect 182791 2931 182839 2959
rect 182529 2897 182839 2931
rect 182529 2869 182577 2897
rect 182605 2869 182639 2897
rect 182667 2869 182701 2897
rect 182729 2869 182763 2897
rect 182791 2869 182839 2897
rect 182529 2835 182839 2869
rect 182529 2807 182577 2835
rect 182605 2807 182639 2835
rect 182667 2807 182701 2835
rect 182729 2807 182763 2835
rect 182791 2807 182839 2835
rect 182529 2773 182839 2807
rect 182529 2745 182577 2773
rect 182605 2745 182639 2773
rect 182667 2745 182701 2773
rect 182729 2745 182763 2773
rect 182791 2745 182839 2773
rect 182529 904 182839 2745
rect 182529 876 182577 904
rect 182605 876 182639 904
rect 182667 876 182701 904
rect 182729 876 182763 904
rect 182791 876 182839 904
rect 182529 842 182839 876
rect 182529 814 182577 842
rect 182605 814 182639 842
rect 182667 814 182701 842
rect 182729 814 182763 842
rect 182791 814 182839 842
rect 182529 780 182839 814
rect 182529 752 182577 780
rect 182605 752 182639 780
rect 182667 752 182701 780
rect 182729 752 182763 780
rect 182791 752 182839 780
rect 182529 718 182839 752
rect 182529 690 182577 718
rect 182605 690 182639 718
rect 182667 690 182701 718
rect 182729 690 182763 718
rect 182791 690 182839 718
rect 182529 162 182839 690
rect 184389 5959 184699 14541
rect 184389 5931 184437 5959
rect 184465 5931 184499 5959
rect 184527 5931 184561 5959
rect 184589 5931 184623 5959
rect 184651 5931 184699 5959
rect 184389 5897 184699 5931
rect 184389 5869 184437 5897
rect 184465 5869 184499 5897
rect 184527 5869 184561 5897
rect 184589 5869 184623 5897
rect 184651 5869 184699 5897
rect 184389 5835 184699 5869
rect 184389 5807 184437 5835
rect 184465 5807 184499 5835
rect 184527 5807 184561 5835
rect 184589 5807 184623 5835
rect 184651 5807 184699 5835
rect 184389 5773 184699 5807
rect 184389 5745 184437 5773
rect 184465 5745 184499 5773
rect 184527 5745 184561 5773
rect 184589 5745 184623 5773
rect 184651 5745 184699 5773
rect 184389 424 184699 5745
rect 184389 396 184437 424
rect 184465 396 184499 424
rect 184527 396 184561 424
rect 184589 396 184623 424
rect 184651 396 184699 424
rect 184389 362 184699 396
rect 184389 334 184437 362
rect 184465 334 184499 362
rect 184527 334 184561 362
rect 184589 334 184623 362
rect 184651 334 184699 362
rect 184389 300 184699 334
rect 184389 272 184437 300
rect 184465 272 184499 300
rect 184527 272 184561 300
rect 184589 272 184623 300
rect 184651 272 184699 300
rect 184389 238 184699 272
rect 184389 210 184437 238
rect 184465 210 184499 238
rect 184527 210 184561 238
rect 184589 210 184623 238
rect 184651 210 184699 238
rect 184389 162 184699 210
rect 191529 11959 191839 14541
rect 191529 11931 191577 11959
rect 191605 11931 191639 11959
rect 191667 11931 191701 11959
rect 191729 11931 191763 11959
rect 191791 11931 191839 11959
rect 191529 11897 191839 11931
rect 191529 11869 191577 11897
rect 191605 11869 191639 11897
rect 191667 11869 191701 11897
rect 191729 11869 191763 11897
rect 191791 11869 191839 11897
rect 191529 11835 191839 11869
rect 191529 11807 191577 11835
rect 191605 11807 191639 11835
rect 191667 11807 191701 11835
rect 191729 11807 191763 11835
rect 191791 11807 191839 11835
rect 191529 11773 191839 11807
rect 191529 11745 191577 11773
rect 191605 11745 191639 11773
rect 191667 11745 191701 11773
rect 191729 11745 191763 11773
rect 191791 11745 191839 11773
rect 191529 2959 191839 11745
rect 191529 2931 191577 2959
rect 191605 2931 191639 2959
rect 191667 2931 191701 2959
rect 191729 2931 191763 2959
rect 191791 2931 191839 2959
rect 191529 2897 191839 2931
rect 191529 2869 191577 2897
rect 191605 2869 191639 2897
rect 191667 2869 191701 2897
rect 191729 2869 191763 2897
rect 191791 2869 191839 2897
rect 191529 2835 191839 2869
rect 191529 2807 191577 2835
rect 191605 2807 191639 2835
rect 191667 2807 191701 2835
rect 191729 2807 191763 2835
rect 191791 2807 191839 2835
rect 191529 2773 191839 2807
rect 191529 2745 191577 2773
rect 191605 2745 191639 2773
rect 191667 2745 191701 2773
rect 191729 2745 191763 2773
rect 191791 2745 191839 2773
rect 191529 904 191839 2745
rect 191529 876 191577 904
rect 191605 876 191639 904
rect 191667 876 191701 904
rect 191729 876 191763 904
rect 191791 876 191839 904
rect 191529 842 191839 876
rect 191529 814 191577 842
rect 191605 814 191639 842
rect 191667 814 191701 842
rect 191729 814 191763 842
rect 191791 814 191839 842
rect 191529 780 191839 814
rect 191529 752 191577 780
rect 191605 752 191639 780
rect 191667 752 191701 780
rect 191729 752 191763 780
rect 191791 752 191839 780
rect 191529 718 191839 752
rect 191529 690 191577 718
rect 191605 690 191639 718
rect 191667 690 191701 718
rect 191729 690 191763 718
rect 191791 690 191839 718
rect 191529 162 191839 690
rect 193389 5959 193699 14541
rect 193389 5931 193437 5959
rect 193465 5931 193499 5959
rect 193527 5931 193561 5959
rect 193589 5931 193623 5959
rect 193651 5931 193699 5959
rect 193389 5897 193699 5931
rect 193389 5869 193437 5897
rect 193465 5869 193499 5897
rect 193527 5869 193561 5897
rect 193589 5869 193623 5897
rect 193651 5869 193699 5897
rect 193389 5835 193699 5869
rect 193389 5807 193437 5835
rect 193465 5807 193499 5835
rect 193527 5807 193561 5835
rect 193589 5807 193623 5835
rect 193651 5807 193699 5835
rect 193389 5773 193699 5807
rect 193389 5745 193437 5773
rect 193465 5745 193499 5773
rect 193527 5745 193561 5773
rect 193589 5745 193623 5773
rect 193651 5745 193699 5773
rect 193389 424 193699 5745
rect 193389 396 193437 424
rect 193465 396 193499 424
rect 193527 396 193561 424
rect 193589 396 193623 424
rect 193651 396 193699 424
rect 193389 362 193699 396
rect 193389 334 193437 362
rect 193465 334 193499 362
rect 193527 334 193561 362
rect 193589 334 193623 362
rect 193651 334 193699 362
rect 193389 300 193699 334
rect 193389 272 193437 300
rect 193465 272 193499 300
rect 193527 272 193561 300
rect 193589 272 193623 300
rect 193651 272 193699 300
rect 193389 238 193699 272
rect 193389 210 193437 238
rect 193465 210 193499 238
rect 193527 210 193561 238
rect 193589 210 193623 238
rect 193651 210 193699 238
rect 193389 162 193699 210
rect 200529 11959 200839 14541
rect 200529 11931 200577 11959
rect 200605 11931 200639 11959
rect 200667 11931 200701 11959
rect 200729 11931 200763 11959
rect 200791 11931 200839 11959
rect 200529 11897 200839 11931
rect 200529 11869 200577 11897
rect 200605 11869 200639 11897
rect 200667 11869 200701 11897
rect 200729 11869 200763 11897
rect 200791 11869 200839 11897
rect 200529 11835 200839 11869
rect 200529 11807 200577 11835
rect 200605 11807 200639 11835
rect 200667 11807 200701 11835
rect 200729 11807 200763 11835
rect 200791 11807 200839 11835
rect 200529 11773 200839 11807
rect 200529 11745 200577 11773
rect 200605 11745 200639 11773
rect 200667 11745 200701 11773
rect 200729 11745 200763 11773
rect 200791 11745 200839 11773
rect 200529 2959 200839 11745
rect 200529 2931 200577 2959
rect 200605 2931 200639 2959
rect 200667 2931 200701 2959
rect 200729 2931 200763 2959
rect 200791 2931 200839 2959
rect 200529 2897 200839 2931
rect 200529 2869 200577 2897
rect 200605 2869 200639 2897
rect 200667 2869 200701 2897
rect 200729 2869 200763 2897
rect 200791 2869 200839 2897
rect 200529 2835 200839 2869
rect 200529 2807 200577 2835
rect 200605 2807 200639 2835
rect 200667 2807 200701 2835
rect 200729 2807 200763 2835
rect 200791 2807 200839 2835
rect 200529 2773 200839 2807
rect 200529 2745 200577 2773
rect 200605 2745 200639 2773
rect 200667 2745 200701 2773
rect 200729 2745 200763 2773
rect 200791 2745 200839 2773
rect 200529 904 200839 2745
rect 200529 876 200577 904
rect 200605 876 200639 904
rect 200667 876 200701 904
rect 200729 876 200763 904
rect 200791 876 200839 904
rect 200529 842 200839 876
rect 200529 814 200577 842
rect 200605 814 200639 842
rect 200667 814 200701 842
rect 200729 814 200763 842
rect 200791 814 200839 842
rect 200529 780 200839 814
rect 200529 752 200577 780
rect 200605 752 200639 780
rect 200667 752 200701 780
rect 200729 752 200763 780
rect 200791 752 200839 780
rect 200529 718 200839 752
rect 200529 690 200577 718
rect 200605 690 200639 718
rect 200667 690 200701 718
rect 200729 690 200763 718
rect 200791 690 200839 718
rect 200529 162 200839 690
rect 202389 5959 202699 14541
rect 202389 5931 202437 5959
rect 202465 5931 202499 5959
rect 202527 5931 202561 5959
rect 202589 5931 202623 5959
rect 202651 5931 202699 5959
rect 202389 5897 202699 5931
rect 202389 5869 202437 5897
rect 202465 5869 202499 5897
rect 202527 5869 202561 5897
rect 202589 5869 202623 5897
rect 202651 5869 202699 5897
rect 202389 5835 202699 5869
rect 202389 5807 202437 5835
rect 202465 5807 202499 5835
rect 202527 5807 202561 5835
rect 202589 5807 202623 5835
rect 202651 5807 202699 5835
rect 202389 5773 202699 5807
rect 202389 5745 202437 5773
rect 202465 5745 202499 5773
rect 202527 5745 202561 5773
rect 202589 5745 202623 5773
rect 202651 5745 202699 5773
rect 202389 424 202699 5745
rect 202389 396 202437 424
rect 202465 396 202499 424
rect 202527 396 202561 424
rect 202589 396 202623 424
rect 202651 396 202699 424
rect 202389 362 202699 396
rect 202389 334 202437 362
rect 202465 334 202499 362
rect 202527 334 202561 362
rect 202589 334 202623 362
rect 202651 334 202699 362
rect 202389 300 202699 334
rect 202389 272 202437 300
rect 202465 272 202499 300
rect 202527 272 202561 300
rect 202589 272 202623 300
rect 202651 272 202699 300
rect 202389 238 202699 272
rect 202389 210 202437 238
rect 202465 210 202499 238
rect 202527 210 202561 238
rect 202589 210 202623 238
rect 202651 210 202699 238
rect 202389 162 202699 210
rect 209529 11959 209839 14541
rect 209529 11931 209577 11959
rect 209605 11931 209639 11959
rect 209667 11931 209701 11959
rect 209729 11931 209763 11959
rect 209791 11931 209839 11959
rect 209529 11897 209839 11931
rect 209529 11869 209577 11897
rect 209605 11869 209639 11897
rect 209667 11869 209701 11897
rect 209729 11869 209763 11897
rect 209791 11869 209839 11897
rect 209529 11835 209839 11869
rect 209529 11807 209577 11835
rect 209605 11807 209639 11835
rect 209667 11807 209701 11835
rect 209729 11807 209763 11835
rect 209791 11807 209839 11835
rect 209529 11773 209839 11807
rect 209529 11745 209577 11773
rect 209605 11745 209639 11773
rect 209667 11745 209701 11773
rect 209729 11745 209763 11773
rect 209791 11745 209839 11773
rect 209529 2959 209839 11745
rect 209529 2931 209577 2959
rect 209605 2931 209639 2959
rect 209667 2931 209701 2959
rect 209729 2931 209763 2959
rect 209791 2931 209839 2959
rect 209529 2897 209839 2931
rect 209529 2869 209577 2897
rect 209605 2869 209639 2897
rect 209667 2869 209701 2897
rect 209729 2869 209763 2897
rect 209791 2869 209839 2897
rect 209529 2835 209839 2869
rect 209529 2807 209577 2835
rect 209605 2807 209639 2835
rect 209667 2807 209701 2835
rect 209729 2807 209763 2835
rect 209791 2807 209839 2835
rect 209529 2773 209839 2807
rect 209529 2745 209577 2773
rect 209605 2745 209639 2773
rect 209667 2745 209701 2773
rect 209729 2745 209763 2773
rect 209791 2745 209839 2773
rect 209529 904 209839 2745
rect 209529 876 209577 904
rect 209605 876 209639 904
rect 209667 876 209701 904
rect 209729 876 209763 904
rect 209791 876 209839 904
rect 209529 842 209839 876
rect 209529 814 209577 842
rect 209605 814 209639 842
rect 209667 814 209701 842
rect 209729 814 209763 842
rect 209791 814 209839 842
rect 209529 780 209839 814
rect 209529 752 209577 780
rect 209605 752 209639 780
rect 209667 752 209701 780
rect 209729 752 209763 780
rect 209791 752 209839 780
rect 209529 718 209839 752
rect 209529 690 209577 718
rect 209605 690 209639 718
rect 209667 690 209701 718
rect 209729 690 209763 718
rect 209791 690 209839 718
rect 209529 162 209839 690
rect 211389 5959 211699 14541
rect 211389 5931 211437 5959
rect 211465 5931 211499 5959
rect 211527 5931 211561 5959
rect 211589 5931 211623 5959
rect 211651 5931 211699 5959
rect 211389 5897 211699 5931
rect 211389 5869 211437 5897
rect 211465 5869 211499 5897
rect 211527 5869 211561 5897
rect 211589 5869 211623 5897
rect 211651 5869 211699 5897
rect 211389 5835 211699 5869
rect 211389 5807 211437 5835
rect 211465 5807 211499 5835
rect 211527 5807 211561 5835
rect 211589 5807 211623 5835
rect 211651 5807 211699 5835
rect 211389 5773 211699 5807
rect 211389 5745 211437 5773
rect 211465 5745 211499 5773
rect 211527 5745 211561 5773
rect 211589 5745 211623 5773
rect 211651 5745 211699 5773
rect 211389 424 211699 5745
rect 211389 396 211437 424
rect 211465 396 211499 424
rect 211527 396 211561 424
rect 211589 396 211623 424
rect 211651 396 211699 424
rect 211389 362 211699 396
rect 211389 334 211437 362
rect 211465 334 211499 362
rect 211527 334 211561 362
rect 211589 334 211623 362
rect 211651 334 211699 362
rect 211389 300 211699 334
rect 211389 272 211437 300
rect 211465 272 211499 300
rect 211527 272 211561 300
rect 211589 272 211623 300
rect 211651 272 211699 300
rect 211389 238 211699 272
rect 211389 210 211437 238
rect 211465 210 211499 238
rect 211527 210 211561 238
rect 211589 210 211623 238
rect 211651 210 211699 238
rect 211389 162 211699 210
rect 218529 11959 218839 14541
rect 218529 11931 218577 11959
rect 218605 11931 218639 11959
rect 218667 11931 218701 11959
rect 218729 11931 218763 11959
rect 218791 11931 218839 11959
rect 218529 11897 218839 11931
rect 218529 11869 218577 11897
rect 218605 11869 218639 11897
rect 218667 11869 218701 11897
rect 218729 11869 218763 11897
rect 218791 11869 218839 11897
rect 218529 11835 218839 11869
rect 218529 11807 218577 11835
rect 218605 11807 218639 11835
rect 218667 11807 218701 11835
rect 218729 11807 218763 11835
rect 218791 11807 218839 11835
rect 218529 11773 218839 11807
rect 218529 11745 218577 11773
rect 218605 11745 218639 11773
rect 218667 11745 218701 11773
rect 218729 11745 218763 11773
rect 218791 11745 218839 11773
rect 218529 2959 218839 11745
rect 218529 2931 218577 2959
rect 218605 2931 218639 2959
rect 218667 2931 218701 2959
rect 218729 2931 218763 2959
rect 218791 2931 218839 2959
rect 218529 2897 218839 2931
rect 218529 2869 218577 2897
rect 218605 2869 218639 2897
rect 218667 2869 218701 2897
rect 218729 2869 218763 2897
rect 218791 2869 218839 2897
rect 218529 2835 218839 2869
rect 218529 2807 218577 2835
rect 218605 2807 218639 2835
rect 218667 2807 218701 2835
rect 218729 2807 218763 2835
rect 218791 2807 218839 2835
rect 218529 2773 218839 2807
rect 218529 2745 218577 2773
rect 218605 2745 218639 2773
rect 218667 2745 218701 2773
rect 218729 2745 218763 2773
rect 218791 2745 218839 2773
rect 218529 904 218839 2745
rect 218529 876 218577 904
rect 218605 876 218639 904
rect 218667 876 218701 904
rect 218729 876 218763 904
rect 218791 876 218839 904
rect 218529 842 218839 876
rect 218529 814 218577 842
rect 218605 814 218639 842
rect 218667 814 218701 842
rect 218729 814 218763 842
rect 218791 814 218839 842
rect 218529 780 218839 814
rect 218529 752 218577 780
rect 218605 752 218639 780
rect 218667 752 218701 780
rect 218729 752 218763 780
rect 218791 752 218839 780
rect 218529 718 218839 752
rect 218529 690 218577 718
rect 218605 690 218639 718
rect 218667 690 218701 718
rect 218729 690 218763 718
rect 218791 690 218839 718
rect 218529 162 218839 690
rect 220389 5959 220699 14541
rect 220389 5931 220437 5959
rect 220465 5931 220499 5959
rect 220527 5931 220561 5959
rect 220589 5931 220623 5959
rect 220651 5931 220699 5959
rect 220389 5897 220699 5931
rect 220389 5869 220437 5897
rect 220465 5869 220499 5897
rect 220527 5869 220561 5897
rect 220589 5869 220623 5897
rect 220651 5869 220699 5897
rect 220389 5835 220699 5869
rect 220389 5807 220437 5835
rect 220465 5807 220499 5835
rect 220527 5807 220561 5835
rect 220589 5807 220623 5835
rect 220651 5807 220699 5835
rect 220389 5773 220699 5807
rect 220389 5745 220437 5773
rect 220465 5745 220499 5773
rect 220527 5745 220561 5773
rect 220589 5745 220623 5773
rect 220651 5745 220699 5773
rect 220389 424 220699 5745
rect 220389 396 220437 424
rect 220465 396 220499 424
rect 220527 396 220561 424
rect 220589 396 220623 424
rect 220651 396 220699 424
rect 220389 362 220699 396
rect 220389 334 220437 362
rect 220465 334 220499 362
rect 220527 334 220561 362
rect 220589 334 220623 362
rect 220651 334 220699 362
rect 220389 300 220699 334
rect 220389 272 220437 300
rect 220465 272 220499 300
rect 220527 272 220561 300
rect 220589 272 220623 300
rect 220651 272 220699 300
rect 220389 238 220699 272
rect 220389 210 220437 238
rect 220465 210 220499 238
rect 220527 210 220561 238
rect 220589 210 220623 238
rect 220651 210 220699 238
rect 220389 162 220699 210
rect 227529 11959 227839 14541
rect 227529 11931 227577 11959
rect 227605 11931 227639 11959
rect 227667 11931 227701 11959
rect 227729 11931 227763 11959
rect 227791 11931 227839 11959
rect 227529 11897 227839 11931
rect 227529 11869 227577 11897
rect 227605 11869 227639 11897
rect 227667 11869 227701 11897
rect 227729 11869 227763 11897
rect 227791 11869 227839 11897
rect 227529 11835 227839 11869
rect 227529 11807 227577 11835
rect 227605 11807 227639 11835
rect 227667 11807 227701 11835
rect 227729 11807 227763 11835
rect 227791 11807 227839 11835
rect 227529 11773 227839 11807
rect 227529 11745 227577 11773
rect 227605 11745 227639 11773
rect 227667 11745 227701 11773
rect 227729 11745 227763 11773
rect 227791 11745 227839 11773
rect 227529 2959 227839 11745
rect 227529 2931 227577 2959
rect 227605 2931 227639 2959
rect 227667 2931 227701 2959
rect 227729 2931 227763 2959
rect 227791 2931 227839 2959
rect 227529 2897 227839 2931
rect 227529 2869 227577 2897
rect 227605 2869 227639 2897
rect 227667 2869 227701 2897
rect 227729 2869 227763 2897
rect 227791 2869 227839 2897
rect 227529 2835 227839 2869
rect 227529 2807 227577 2835
rect 227605 2807 227639 2835
rect 227667 2807 227701 2835
rect 227729 2807 227763 2835
rect 227791 2807 227839 2835
rect 227529 2773 227839 2807
rect 227529 2745 227577 2773
rect 227605 2745 227639 2773
rect 227667 2745 227701 2773
rect 227729 2745 227763 2773
rect 227791 2745 227839 2773
rect 227529 904 227839 2745
rect 227529 876 227577 904
rect 227605 876 227639 904
rect 227667 876 227701 904
rect 227729 876 227763 904
rect 227791 876 227839 904
rect 227529 842 227839 876
rect 227529 814 227577 842
rect 227605 814 227639 842
rect 227667 814 227701 842
rect 227729 814 227763 842
rect 227791 814 227839 842
rect 227529 780 227839 814
rect 227529 752 227577 780
rect 227605 752 227639 780
rect 227667 752 227701 780
rect 227729 752 227763 780
rect 227791 752 227839 780
rect 227529 718 227839 752
rect 227529 690 227577 718
rect 227605 690 227639 718
rect 227667 690 227701 718
rect 227729 690 227763 718
rect 227791 690 227839 718
rect 227529 162 227839 690
rect 229389 5959 229699 14541
rect 229389 5931 229437 5959
rect 229465 5931 229499 5959
rect 229527 5931 229561 5959
rect 229589 5931 229623 5959
rect 229651 5931 229699 5959
rect 229389 5897 229699 5931
rect 229389 5869 229437 5897
rect 229465 5869 229499 5897
rect 229527 5869 229561 5897
rect 229589 5869 229623 5897
rect 229651 5869 229699 5897
rect 229389 5835 229699 5869
rect 229389 5807 229437 5835
rect 229465 5807 229499 5835
rect 229527 5807 229561 5835
rect 229589 5807 229623 5835
rect 229651 5807 229699 5835
rect 229389 5773 229699 5807
rect 229389 5745 229437 5773
rect 229465 5745 229499 5773
rect 229527 5745 229561 5773
rect 229589 5745 229623 5773
rect 229651 5745 229699 5773
rect 229389 424 229699 5745
rect 229389 396 229437 424
rect 229465 396 229499 424
rect 229527 396 229561 424
rect 229589 396 229623 424
rect 229651 396 229699 424
rect 229389 362 229699 396
rect 229389 334 229437 362
rect 229465 334 229499 362
rect 229527 334 229561 362
rect 229589 334 229623 362
rect 229651 334 229699 362
rect 229389 300 229699 334
rect 229389 272 229437 300
rect 229465 272 229499 300
rect 229527 272 229561 300
rect 229589 272 229623 300
rect 229651 272 229699 300
rect 229389 238 229699 272
rect 229389 210 229437 238
rect 229465 210 229499 238
rect 229527 210 229561 238
rect 229589 210 229623 238
rect 229651 210 229699 238
rect 229389 162 229699 210
rect 236529 11959 236839 14541
rect 236529 11931 236577 11959
rect 236605 11931 236639 11959
rect 236667 11931 236701 11959
rect 236729 11931 236763 11959
rect 236791 11931 236839 11959
rect 236529 11897 236839 11931
rect 236529 11869 236577 11897
rect 236605 11869 236639 11897
rect 236667 11869 236701 11897
rect 236729 11869 236763 11897
rect 236791 11869 236839 11897
rect 236529 11835 236839 11869
rect 236529 11807 236577 11835
rect 236605 11807 236639 11835
rect 236667 11807 236701 11835
rect 236729 11807 236763 11835
rect 236791 11807 236839 11835
rect 236529 11773 236839 11807
rect 236529 11745 236577 11773
rect 236605 11745 236639 11773
rect 236667 11745 236701 11773
rect 236729 11745 236763 11773
rect 236791 11745 236839 11773
rect 236529 2959 236839 11745
rect 236529 2931 236577 2959
rect 236605 2931 236639 2959
rect 236667 2931 236701 2959
rect 236729 2931 236763 2959
rect 236791 2931 236839 2959
rect 236529 2897 236839 2931
rect 236529 2869 236577 2897
rect 236605 2869 236639 2897
rect 236667 2869 236701 2897
rect 236729 2869 236763 2897
rect 236791 2869 236839 2897
rect 236529 2835 236839 2869
rect 236529 2807 236577 2835
rect 236605 2807 236639 2835
rect 236667 2807 236701 2835
rect 236729 2807 236763 2835
rect 236791 2807 236839 2835
rect 236529 2773 236839 2807
rect 236529 2745 236577 2773
rect 236605 2745 236639 2773
rect 236667 2745 236701 2773
rect 236729 2745 236763 2773
rect 236791 2745 236839 2773
rect 236529 904 236839 2745
rect 236529 876 236577 904
rect 236605 876 236639 904
rect 236667 876 236701 904
rect 236729 876 236763 904
rect 236791 876 236839 904
rect 236529 842 236839 876
rect 236529 814 236577 842
rect 236605 814 236639 842
rect 236667 814 236701 842
rect 236729 814 236763 842
rect 236791 814 236839 842
rect 236529 780 236839 814
rect 236529 752 236577 780
rect 236605 752 236639 780
rect 236667 752 236701 780
rect 236729 752 236763 780
rect 236791 752 236839 780
rect 236529 718 236839 752
rect 236529 690 236577 718
rect 236605 690 236639 718
rect 236667 690 236701 718
rect 236729 690 236763 718
rect 236791 690 236839 718
rect 236529 162 236839 690
rect 238389 5959 238699 14541
rect 238389 5931 238437 5959
rect 238465 5931 238499 5959
rect 238527 5931 238561 5959
rect 238589 5931 238623 5959
rect 238651 5931 238699 5959
rect 238389 5897 238699 5931
rect 238389 5869 238437 5897
rect 238465 5869 238499 5897
rect 238527 5869 238561 5897
rect 238589 5869 238623 5897
rect 238651 5869 238699 5897
rect 238389 5835 238699 5869
rect 238389 5807 238437 5835
rect 238465 5807 238499 5835
rect 238527 5807 238561 5835
rect 238589 5807 238623 5835
rect 238651 5807 238699 5835
rect 238389 5773 238699 5807
rect 238389 5745 238437 5773
rect 238465 5745 238499 5773
rect 238527 5745 238561 5773
rect 238589 5745 238623 5773
rect 238651 5745 238699 5773
rect 238389 424 238699 5745
rect 238389 396 238437 424
rect 238465 396 238499 424
rect 238527 396 238561 424
rect 238589 396 238623 424
rect 238651 396 238699 424
rect 238389 362 238699 396
rect 238389 334 238437 362
rect 238465 334 238499 362
rect 238527 334 238561 362
rect 238589 334 238623 362
rect 238651 334 238699 362
rect 238389 300 238699 334
rect 238389 272 238437 300
rect 238465 272 238499 300
rect 238527 272 238561 300
rect 238589 272 238623 300
rect 238651 272 238699 300
rect 238389 238 238699 272
rect 238389 210 238437 238
rect 238465 210 238499 238
rect 238527 210 238561 238
rect 238589 210 238623 238
rect 238651 210 238699 238
rect 238389 162 238699 210
rect 245529 11959 245839 14541
rect 245529 11931 245577 11959
rect 245605 11931 245639 11959
rect 245667 11931 245701 11959
rect 245729 11931 245763 11959
rect 245791 11931 245839 11959
rect 245529 11897 245839 11931
rect 245529 11869 245577 11897
rect 245605 11869 245639 11897
rect 245667 11869 245701 11897
rect 245729 11869 245763 11897
rect 245791 11869 245839 11897
rect 245529 11835 245839 11869
rect 245529 11807 245577 11835
rect 245605 11807 245639 11835
rect 245667 11807 245701 11835
rect 245729 11807 245763 11835
rect 245791 11807 245839 11835
rect 245529 11773 245839 11807
rect 245529 11745 245577 11773
rect 245605 11745 245639 11773
rect 245667 11745 245701 11773
rect 245729 11745 245763 11773
rect 245791 11745 245839 11773
rect 245529 2959 245839 11745
rect 245529 2931 245577 2959
rect 245605 2931 245639 2959
rect 245667 2931 245701 2959
rect 245729 2931 245763 2959
rect 245791 2931 245839 2959
rect 245529 2897 245839 2931
rect 245529 2869 245577 2897
rect 245605 2869 245639 2897
rect 245667 2869 245701 2897
rect 245729 2869 245763 2897
rect 245791 2869 245839 2897
rect 245529 2835 245839 2869
rect 245529 2807 245577 2835
rect 245605 2807 245639 2835
rect 245667 2807 245701 2835
rect 245729 2807 245763 2835
rect 245791 2807 245839 2835
rect 245529 2773 245839 2807
rect 245529 2745 245577 2773
rect 245605 2745 245639 2773
rect 245667 2745 245701 2773
rect 245729 2745 245763 2773
rect 245791 2745 245839 2773
rect 245529 904 245839 2745
rect 245529 876 245577 904
rect 245605 876 245639 904
rect 245667 876 245701 904
rect 245729 876 245763 904
rect 245791 876 245839 904
rect 245529 842 245839 876
rect 245529 814 245577 842
rect 245605 814 245639 842
rect 245667 814 245701 842
rect 245729 814 245763 842
rect 245791 814 245839 842
rect 245529 780 245839 814
rect 245529 752 245577 780
rect 245605 752 245639 780
rect 245667 752 245701 780
rect 245729 752 245763 780
rect 245791 752 245839 780
rect 245529 718 245839 752
rect 245529 690 245577 718
rect 245605 690 245639 718
rect 245667 690 245701 718
rect 245729 690 245763 718
rect 245791 690 245839 718
rect 245529 162 245839 690
rect 247389 5959 247699 14745
rect 247389 5931 247437 5959
rect 247465 5931 247499 5959
rect 247527 5931 247561 5959
rect 247589 5931 247623 5959
rect 247651 5931 247699 5959
rect 247389 5897 247699 5931
rect 247389 5869 247437 5897
rect 247465 5869 247499 5897
rect 247527 5869 247561 5897
rect 247589 5869 247623 5897
rect 247651 5869 247699 5897
rect 247389 5835 247699 5869
rect 247389 5807 247437 5835
rect 247465 5807 247499 5835
rect 247527 5807 247561 5835
rect 247589 5807 247623 5835
rect 247651 5807 247699 5835
rect 247389 5773 247699 5807
rect 247389 5745 247437 5773
rect 247465 5745 247499 5773
rect 247527 5745 247561 5773
rect 247589 5745 247623 5773
rect 247651 5745 247699 5773
rect 247389 424 247699 5745
rect 247389 396 247437 424
rect 247465 396 247499 424
rect 247527 396 247561 424
rect 247589 396 247623 424
rect 247651 396 247699 424
rect 247389 362 247699 396
rect 247389 334 247437 362
rect 247465 334 247499 362
rect 247527 334 247561 362
rect 247589 334 247623 362
rect 247651 334 247699 362
rect 247389 300 247699 334
rect 247389 272 247437 300
rect 247465 272 247499 300
rect 247527 272 247561 300
rect 247589 272 247623 300
rect 247651 272 247699 300
rect 247389 238 247699 272
rect 247389 210 247437 238
rect 247465 210 247499 238
rect 247527 210 247561 238
rect 247589 210 247623 238
rect 247651 210 247699 238
rect 247389 162 247699 210
rect 254529 11959 254839 20745
rect 254870 256634 254898 256639
rect 254870 14210 254898 256606
rect 254870 14177 254898 14182
rect 256389 248959 256699 257745
rect 256389 248931 256437 248959
rect 256465 248931 256499 248959
rect 256527 248931 256561 248959
rect 256589 248931 256623 248959
rect 256651 248931 256699 248959
rect 256389 248897 256699 248931
rect 256389 248869 256437 248897
rect 256465 248869 256499 248897
rect 256527 248869 256561 248897
rect 256589 248869 256623 248897
rect 256651 248869 256699 248897
rect 256389 248835 256699 248869
rect 256389 248807 256437 248835
rect 256465 248807 256499 248835
rect 256527 248807 256561 248835
rect 256589 248807 256623 248835
rect 256651 248807 256699 248835
rect 256389 248773 256699 248807
rect 256389 248745 256437 248773
rect 256465 248745 256499 248773
rect 256527 248745 256561 248773
rect 256589 248745 256623 248773
rect 256651 248745 256699 248773
rect 256389 239959 256699 248745
rect 256389 239931 256437 239959
rect 256465 239931 256499 239959
rect 256527 239931 256561 239959
rect 256589 239931 256623 239959
rect 256651 239931 256699 239959
rect 256389 239897 256699 239931
rect 256389 239869 256437 239897
rect 256465 239869 256499 239897
rect 256527 239869 256561 239897
rect 256589 239869 256623 239897
rect 256651 239869 256699 239897
rect 256389 239835 256699 239869
rect 256389 239807 256437 239835
rect 256465 239807 256499 239835
rect 256527 239807 256561 239835
rect 256589 239807 256623 239835
rect 256651 239807 256699 239835
rect 256389 239773 256699 239807
rect 256389 239745 256437 239773
rect 256465 239745 256499 239773
rect 256527 239745 256561 239773
rect 256589 239745 256623 239773
rect 256651 239745 256699 239773
rect 256389 230959 256699 239745
rect 256389 230931 256437 230959
rect 256465 230931 256499 230959
rect 256527 230931 256561 230959
rect 256589 230931 256623 230959
rect 256651 230931 256699 230959
rect 256389 230897 256699 230931
rect 256389 230869 256437 230897
rect 256465 230869 256499 230897
rect 256527 230869 256561 230897
rect 256589 230869 256623 230897
rect 256651 230869 256699 230897
rect 256389 230835 256699 230869
rect 256389 230807 256437 230835
rect 256465 230807 256499 230835
rect 256527 230807 256561 230835
rect 256589 230807 256623 230835
rect 256651 230807 256699 230835
rect 256389 230773 256699 230807
rect 256389 230745 256437 230773
rect 256465 230745 256499 230773
rect 256527 230745 256561 230773
rect 256589 230745 256623 230773
rect 256651 230745 256699 230773
rect 256389 221959 256699 230745
rect 256389 221931 256437 221959
rect 256465 221931 256499 221959
rect 256527 221931 256561 221959
rect 256589 221931 256623 221959
rect 256651 221931 256699 221959
rect 256389 221897 256699 221931
rect 256389 221869 256437 221897
rect 256465 221869 256499 221897
rect 256527 221869 256561 221897
rect 256589 221869 256623 221897
rect 256651 221869 256699 221897
rect 256389 221835 256699 221869
rect 256389 221807 256437 221835
rect 256465 221807 256499 221835
rect 256527 221807 256561 221835
rect 256589 221807 256623 221835
rect 256651 221807 256699 221835
rect 256389 221773 256699 221807
rect 256389 221745 256437 221773
rect 256465 221745 256499 221773
rect 256527 221745 256561 221773
rect 256589 221745 256623 221773
rect 256651 221745 256699 221773
rect 256389 212959 256699 221745
rect 256389 212931 256437 212959
rect 256465 212931 256499 212959
rect 256527 212931 256561 212959
rect 256589 212931 256623 212959
rect 256651 212931 256699 212959
rect 256389 212897 256699 212931
rect 256389 212869 256437 212897
rect 256465 212869 256499 212897
rect 256527 212869 256561 212897
rect 256589 212869 256623 212897
rect 256651 212869 256699 212897
rect 256389 212835 256699 212869
rect 256389 212807 256437 212835
rect 256465 212807 256499 212835
rect 256527 212807 256561 212835
rect 256589 212807 256623 212835
rect 256651 212807 256699 212835
rect 256389 212773 256699 212807
rect 256389 212745 256437 212773
rect 256465 212745 256499 212773
rect 256527 212745 256561 212773
rect 256589 212745 256623 212773
rect 256651 212745 256699 212773
rect 256389 203959 256699 212745
rect 256389 203931 256437 203959
rect 256465 203931 256499 203959
rect 256527 203931 256561 203959
rect 256589 203931 256623 203959
rect 256651 203931 256699 203959
rect 256389 203897 256699 203931
rect 256389 203869 256437 203897
rect 256465 203869 256499 203897
rect 256527 203869 256561 203897
rect 256589 203869 256623 203897
rect 256651 203869 256699 203897
rect 256389 203835 256699 203869
rect 256389 203807 256437 203835
rect 256465 203807 256499 203835
rect 256527 203807 256561 203835
rect 256589 203807 256623 203835
rect 256651 203807 256699 203835
rect 256389 203773 256699 203807
rect 256389 203745 256437 203773
rect 256465 203745 256499 203773
rect 256527 203745 256561 203773
rect 256589 203745 256623 203773
rect 256651 203745 256699 203773
rect 256389 194959 256699 203745
rect 256389 194931 256437 194959
rect 256465 194931 256499 194959
rect 256527 194931 256561 194959
rect 256589 194931 256623 194959
rect 256651 194931 256699 194959
rect 256389 194897 256699 194931
rect 256389 194869 256437 194897
rect 256465 194869 256499 194897
rect 256527 194869 256561 194897
rect 256589 194869 256623 194897
rect 256651 194869 256699 194897
rect 256389 194835 256699 194869
rect 256389 194807 256437 194835
rect 256465 194807 256499 194835
rect 256527 194807 256561 194835
rect 256589 194807 256623 194835
rect 256651 194807 256699 194835
rect 256389 194773 256699 194807
rect 256389 194745 256437 194773
rect 256465 194745 256499 194773
rect 256527 194745 256561 194773
rect 256589 194745 256623 194773
rect 256651 194745 256699 194773
rect 256389 185959 256699 194745
rect 256389 185931 256437 185959
rect 256465 185931 256499 185959
rect 256527 185931 256561 185959
rect 256589 185931 256623 185959
rect 256651 185931 256699 185959
rect 256389 185897 256699 185931
rect 256389 185869 256437 185897
rect 256465 185869 256499 185897
rect 256527 185869 256561 185897
rect 256589 185869 256623 185897
rect 256651 185869 256699 185897
rect 256389 185835 256699 185869
rect 256389 185807 256437 185835
rect 256465 185807 256499 185835
rect 256527 185807 256561 185835
rect 256589 185807 256623 185835
rect 256651 185807 256699 185835
rect 256389 185773 256699 185807
rect 256389 185745 256437 185773
rect 256465 185745 256499 185773
rect 256527 185745 256561 185773
rect 256589 185745 256623 185773
rect 256651 185745 256699 185773
rect 256389 176959 256699 185745
rect 256389 176931 256437 176959
rect 256465 176931 256499 176959
rect 256527 176931 256561 176959
rect 256589 176931 256623 176959
rect 256651 176931 256699 176959
rect 256389 176897 256699 176931
rect 256389 176869 256437 176897
rect 256465 176869 256499 176897
rect 256527 176869 256561 176897
rect 256589 176869 256623 176897
rect 256651 176869 256699 176897
rect 256389 176835 256699 176869
rect 256389 176807 256437 176835
rect 256465 176807 256499 176835
rect 256527 176807 256561 176835
rect 256589 176807 256623 176835
rect 256651 176807 256699 176835
rect 256389 176773 256699 176807
rect 256389 176745 256437 176773
rect 256465 176745 256499 176773
rect 256527 176745 256561 176773
rect 256589 176745 256623 176773
rect 256651 176745 256699 176773
rect 256389 167959 256699 176745
rect 256389 167931 256437 167959
rect 256465 167931 256499 167959
rect 256527 167931 256561 167959
rect 256589 167931 256623 167959
rect 256651 167931 256699 167959
rect 256389 167897 256699 167931
rect 256389 167869 256437 167897
rect 256465 167869 256499 167897
rect 256527 167869 256561 167897
rect 256589 167869 256623 167897
rect 256651 167869 256699 167897
rect 256389 167835 256699 167869
rect 256389 167807 256437 167835
rect 256465 167807 256499 167835
rect 256527 167807 256561 167835
rect 256589 167807 256623 167835
rect 256651 167807 256699 167835
rect 256389 167773 256699 167807
rect 256389 167745 256437 167773
rect 256465 167745 256499 167773
rect 256527 167745 256561 167773
rect 256589 167745 256623 167773
rect 256651 167745 256699 167773
rect 256389 158959 256699 167745
rect 256389 158931 256437 158959
rect 256465 158931 256499 158959
rect 256527 158931 256561 158959
rect 256589 158931 256623 158959
rect 256651 158931 256699 158959
rect 256389 158897 256699 158931
rect 256389 158869 256437 158897
rect 256465 158869 256499 158897
rect 256527 158869 256561 158897
rect 256589 158869 256623 158897
rect 256651 158869 256699 158897
rect 256389 158835 256699 158869
rect 256389 158807 256437 158835
rect 256465 158807 256499 158835
rect 256527 158807 256561 158835
rect 256589 158807 256623 158835
rect 256651 158807 256699 158835
rect 256389 158773 256699 158807
rect 256389 158745 256437 158773
rect 256465 158745 256499 158773
rect 256527 158745 256561 158773
rect 256589 158745 256623 158773
rect 256651 158745 256699 158773
rect 256389 149959 256699 158745
rect 256389 149931 256437 149959
rect 256465 149931 256499 149959
rect 256527 149931 256561 149959
rect 256589 149931 256623 149959
rect 256651 149931 256699 149959
rect 256389 149897 256699 149931
rect 256389 149869 256437 149897
rect 256465 149869 256499 149897
rect 256527 149869 256561 149897
rect 256589 149869 256623 149897
rect 256651 149869 256699 149897
rect 256389 149835 256699 149869
rect 256389 149807 256437 149835
rect 256465 149807 256499 149835
rect 256527 149807 256561 149835
rect 256589 149807 256623 149835
rect 256651 149807 256699 149835
rect 256389 149773 256699 149807
rect 256389 149745 256437 149773
rect 256465 149745 256499 149773
rect 256527 149745 256561 149773
rect 256589 149745 256623 149773
rect 256651 149745 256699 149773
rect 256389 140959 256699 149745
rect 256389 140931 256437 140959
rect 256465 140931 256499 140959
rect 256527 140931 256561 140959
rect 256589 140931 256623 140959
rect 256651 140931 256699 140959
rect 256389 140897 256699 140931
rect 256389 140869 256437 140897
rect 256465 140869 256499 140897
rect 256527 140869 256561 140897
rect 256589 140869 256623 140897
rect 256651 140869 256699 140897
rect 256389 140835 256699 140869
rect 256389 140807 256437 140835
rect 256465 140807 256499 140835
rect 256527 140807 256561 140835
rect 256589 140807 256623 140835
rect 256651 140807 256699 140835
rect 256389 140773 256699 140807
rect 256389 140745 256437 140773
rect 256465 140745 256499 140773
rect 256527 140745 256561 140773
rect 256589 140745 256623 140773
rect 256651 140745 256699 140773
rect 256389 131959 256699 140745
rect 256389 131931 256437 131959
rect 256465 131931 256499 131959
rect 256527 131931 256561 131959
rect 256589 131931 256623 131959
rect 256651 131931 256699 131959
rect 256389 131897 256699 131931
rect 256389 131869 256437 131897
rect 256465 131869 256499 131897
rect 256527 131869 256561 131897
rect 256589 131869 256623 131897
rect 256651 131869 256699 131897
rect 256389 131835 256699 131869
rect 256389 131807 256437 131835
rect 256465 131807 256499 131835
rect 256527 131807 256561 131835
rect 256589 131807 256623 131835
rect 256651 131807 256699 131835
rect 256389 131773 256699 131807
rect 256389 131745 256437 131773
rect 256465 131745 256499 131773
rect 256527 131745 256561 131773
rect 256589 131745 256623 131773
rect 256651 131745 256699 131773
rect 256389 122959 256699 131745
rect 256389 122931 256437 122959
rect 256465 122931 256499 122959
rect 256527 122931 256561 122959
rect 256589 122931 256623 122959
rect 256651 122931 256699 122959
rect 256389 122897 256699 122931
rect 256389 122869 256437 122897
rect 256465 122869 256499 122897
rect 256527 122869 256561 122897
rect 256589 122869 256623 122897
rect 256651 122869 256699 122897
rect 256389 122835 256699 122869
rect 256389 122807 256437 122835
rect 256465 122807 256499 122835
rect 256527 122807 256561 122835
rect 256589 122807 256623 122835
rect 256651 122807 256699 122835
rect 256389 122773 256699 122807
rect 256389 122745 256437 122773
rect 256465 122745 256499 122773
rect 256527 122745 256561 122773
rect 256589 122745 256623 122773
rect 256651 122745 256699 122773
rect 256389 113959 256699 122745
rect 256389 113931 256437 113959
rect 256465 113931 256499 113959
rect 256527 113931 256561 113959
rect 256589 113931 256623 113959
rect 256651 113931 256699 113959
rect 256389 113897 256699 113931
rect 256389 113869 256437 113897
rect 256465 113869 256499 113897
rect 256527 113869 256561 113897
rect 256589 113869 256623 113897
rect 256651 113869 256699 113897
rect 256389 113835 256699 113869
rect 256389 113807 256437 113835
rect 256465 113807 256499 113835
rect 256527 113807 256561 113835
rect 256589 113807 256623 113835
rect 256651 113807 256699 113835
rect 256389 113773 256699 113807
rect 256389 113745 256437 113773
rect 256465 113745 256499 113773
rect 256527 113745 256561 113773
rect 256589 113745 256623 113773
rect 256651 113745 256699 113773
rect 256389 104959 256699 113745
rect 256389 104931 256437 104959
rect 256465 104931 256499 104959
rect 256527 104931 256561 104959
rect 256589 104931 256623 104959
rect 256651 104931 256699 104959
rect 256389 104897 256699 104931
rect 256389 104869 256437 104897
rect 256465 104869 256499 104897
rect 256527 104869 256561 104897
rect 256589 104869 256623 104897
rect 256651 104869 256699 104897
rect 256389 104835 256699 104869
rect 256389 104807 256437 104835
rect 256465 104807 256499 104835
rect 256527 104807 256561 104835
rect 256589 104807 256623 104835
rect 256651 104807 256699 104835
rect 256389 104773 256699 104807
rect 256389 104745 256437 104773
rect 256465 104745 256499 104773
rect 256527 104745 256561 104773
rect 256589 104745 256623 104773
rect 256651 104745 256699 104773
rect 256389 95959 256699 104745
rect 256389 95931 256437 95959
rect 256465 95931 256499 95959
rect 256527 95931 256561 95959
rect 256589 95931 256623 95959
rect 256651 95931 256699 95959
rect 256389 95897 256699 95931
rect 256389 95869 256437 95897
rect 256465 95869 256499 95897
rect 256527 95869 256561 95897
rect 256589 95869 256623 95897
rect 256651 95869 256699 95897
rect 256389 95835 256699 95869
rect 256389 95807 256437 95835
rect 256465 95807 256499 95835
rect 256527 95807 256561 95835
rect 256589 95807 256623 95835
rect 256651 95807 256699 95835
rect 256389 95773 256699 95807
rect 256389 95745 256437 95773
rect 256465 95745 256499 95773
rect 256527 95745 256561 95773
rect 256589 95745 256623 95773
rect 256651 95745 256699 95773
rect 256389 86959 256699 95745
rect 256389 86931 256437 86959
rect 256465 86931 256499 86959
rect 256527 86931 256561 86959
rect 256589 86931 256623 86959
rect 256651 86931 256699 86959
rect 256389 86897 256699 86931
rect 256389 86869 256437 86897
rect 256465 86869 256499 86897
rect 256527 86869 256561 86897
rect 256589 86869 256623 86897
rect 256651 86869 256699 86897
rect 256389 86835 256699 86869
rect 256389 86807 256437 86835
rect 256465 86807 256499 86835
rect 256527 86807 256561 86835
rect 256589 86807 256623 86835
rect 256651 86807 256699 86835
rect 256389 86773 256699 86807
rect 256389 86745 256437 86773
rect 256465 86745 256499 86773
rect 256527 86745 256561 86773
rect 256589 86745 256623 86773
rect 256651 86745 256699 86773
rect 256389 77959 256699 86745
rect 256389 77931 256437 77959
rect 256465 77931 256499 77959
rect 256527 77931 256561 77959
rect 256589 77931 256623 77959
rect 256651 77931 256699 77959
rect 256389 77897 256699 77931
rect 256389 77869 256437 77897
rect 256465 77869 256499 77897
rect 256527 77869 256561 77897
rect 256589 77869 256623 77897
rect 256651 77869 256699 77897
rect 256389 77835 256699 77869
rect 256389 77807 256437 77835
rect 256465 77807 256499 77835
rect 256527 77807 256561 77835
rect 256589 77807 256623 77835
rect 256651 77807 256699 77835
rect 256389 77773 256699 77807
rect 256389 77745 256437 77773
rect 256465 77745 256499 77773
rect 256527 77745 256561 77773
rect 256589 77745 256623 77773
rect 256651 77745 256699 77773
rect 256389 68959 256699 77745
rect 256389 68931 256437 68959
rect 256465 68931 256499 68959
rect 256527 68931 256561 68959
rect 256589 68931 256623 68959
rect 256651 68931 256699 68959
rect 256389 68897 256699 68931
rect 256389 68869 256437 68897
rect 256465 68869 256499 68897
rect 256527 68869 256561 68897
rect 256589 68869 256623 68897
rect 256651 68869 256699 68897
rect 256389 68835 256699 68869
rect 256389 68807 256437 68835
rect 256465 68807 256499 68835
rect 256527 68807 256561 68835
rect 256589 68807 256623 68835
rect 256651 68807 256699 68835
rect 256389 68773 256699 68807
rect 256389 68745 256437 68773
rect 256465 68745 256499 68773
rect 256527 68745 256561 68773
rect 256589 68745 256623 68773
rect 256651 68745 256699 68773
rect 256389 59959 256699 68745
rect 256389 59931 256437 59959
rect 256465 59931 256499 59959
rect 256527 59931 256561 59959
rect 256589 59931 256623 59959
rect 256651 59931 256699 59959
rect 256389 59897 256699 59931
rect 256389 59869 256437 59897
rect 256465 59869 256499 59897
rect 256527 59869 256561 59897
rect 256589 59869 256623 59897
rect 256651 59869 256699 59897
rect 256389 59835 256699 59869
rect 256389 59807 256437 59835
rect 256465 59807 256499 59835
rect 256527 59807 256561 59835
rect 256589 59807 256623 59835
rect 256651 59807 256699 59835
rect 256389 59773 256699 59807
rect 256389 59745 256437 59773
rect 256465 59745 256499 59773
rect 256527 59745 256561 59773
rect 256589 59745 256623 59773
rect 256651 59745 256699 59773
rect 256389 50959 256699 59745
rect 256389 50931 256437 50959
rect 256465 50931 256499 50959
rect 256527 50931 256561 50959
rect 256589 50931 256623 50959
rect 256651 50931 256699 50959
rect 256389 50897 256699 50931
rect 256389 50869 256437 50897
rect 256465 50869 256499 50897
rect 256527 50869 256561 50897
rect 256589 50869 256623 50897
rect 256651 50869 256699 50897
rect 256389 50835 256699 50869
rect 256389 50807 256437 50835
rect 256465 50807 256499 50835
rect 256527 50807 256561 50835
rect 256589 50807 256623 50835
rect 256651 50807 256699 50835
rect 256389 50773 256699 50807
rect 256389 50745 256437 50773
rect 256465 50745 256499 50773
rect 256527 50745 256561 50773
rect 256589 50745 256623 50773
rect 256651 50745 256699 50773
rect 256389 41959 256699 50745
rect 256389 41931 256437 41959
rect 256465 41931 256499 41959
rect 256527 41931 256561 41959
rect 256589 41931 256623 41959
rect 256651 41931 256699 41959
rect 256389 41897 256699 41931
rect 256389 41869 256437 41897
rect 256465 41869 256499 41897
rect 256527 41869 256561 41897
rect 256589 41869 256623 41897
rect 256651 41869 256699 41897
rect 256389 41835 256699 41869
rect 256389 41807 256437 41835
rect 256465 41807 256499 41835
rect 256527 41807 256561 41835
rect 256589 41807 256623 41835
rect 256651 41807 256699 41835
rect 256389 41773 256699 41807
rect 256389 41745 256437 41773
rect 256465 41745 256499 41773
rect 256527 41745 256561 41773
rect 256589 41745 256623 41773
rect 256651 41745 256699 41773
rect 256389 32959 256699 41745
rect 256389 32931 256437 32959
rect 256465 32931 256499 32959
rect 256527 32931 256561 32959
rect 256589 32931 256623 32959
rect 256651 32931 256699 32959
rect 256389 32897 256699 32931
rect 256389 32869 256437 32897
rect 256465 32869 256499 32897
rect 256527 32869 256561 32897
rect 256589 32869 256623 32897
rect 256651 32869 256699 32897
rect 256389 32835 256699 32869
rect 256389 32807 256437 32835
rect 256465 32807 256499 32835
rect 256527 32807 256561 32835
rect 256589 32807 256623 32835
rect 256651 32807 256699 32835
rect 256389 32773 256699 32807
rect 256389 32745 256437 32773
rect 256465 32745 256499 32773
rect 256527 32745 256561 32773
rect 256589 32745 256623 32773
rect 256651 32745 256699 32773
rect 256389 23959 256699 32745
rect 256389 23931 256437 23959
rect 256465 23931 256499 23959
rect 256527 23931 256561 23959
rect 256589 23931 256623 23959
rect 256651 23931 256699 23959
rect 256389 23897 256699 23931
rect 256389 23869 256437 23897
rect 256465 23869 256499 23897
rect 256527 23869 256561 23897
rect 256589 23869 256623 23897
rect 256651 23869 256699 23897
rect 256389 23835 256699 23869
rect 256389 23807 256437 23835
rect 256465 23807 256499 23835
rect 256527 23807 256561 23835
rect 256589 23807 256623 23835
rect 256651 23807 256699 23835
rect 256389 23773 256699 23807
rect 256389 23745 256437 23773
rect 256465 23745 256499 23773
rect 256527 23745 256561 23773
rect 256589 23745 256623 23773
rect 256651 23745 256699 23773
rect 256389 14959 256699 23745
rect 256389 14931 256437 14959
rect 256465 14931 256499 14959
rect 256527 14931 256561 14959
rect 256589 14931 256623 14959
rect 256651 14931 256699 14959
rect 256389 14897 256699 14931
rect 256389 14869 256437 14897
rect 256465 14869 256499 14897
rect 256527 14869 256561 14897
rect 256589 14869 256623 14897
rect 256651 14869 256699 14897
rect 256389 14835 256699 14869
rect 256389 14807 256437 14835
rect 256465 14807 256499 14835
rect 256527 14807 256561 14835
rect 256589 14807 256623 14835
rect 256651 14807 256699 14835
rect 256389 14773 256699 14807
rect 256389 14745 256437 14773
rect 256465 14745 256499 14773
rect 256527 14745 256561 14773
rect 256589 14745 256623 14773
rect 256651 14745 256699 14773
rect 254529 11931 254577 11959
rect 254605 11931 254639 11959
rect 254667 11931 254701 11959
rect 254729 11931 254763 11959
rect 254791 11931 254839 11959
rect 254529 11897 254839 11931
rect 254529 11869 254577 11897
rect 254605 11869 254639 11897
rect 254667 11869 254701 11897
rect 254729 11869 254763 11897
rect 254791 11869 254839 11897
rect 254529 11835 254839 11869
rect 254529 11807 254577 11835
rect 254605 11807 254639 11835
rect 254667 11807 254701 11835
rect 254729 11807 254763 11835
rect 254791 11807 254839 11835
rect 254529 11773 254839 11807
rect 254529 11745 254577 11773
rect 254605 11745 254639 11773
rect 254667 11745 254701 11773
rect 254729 11745 254763 11773
rect 254791 11745 254839 11773
rect 254529 2959 254839 11745
rect 254529 2931 254577 2959
rect 254605 2931 254639 2959
rect 254667 2931 254701 2959
rect 254729 2931 254763 2959
rect 254791 2931 254839 2959
rect 254529 2897 254839 2931
rect 254529 2869 254577 2897
rect 254605 2869 254639 2897
rect 254667 2869 254701 2897
rect 254729 2869 254763 2897
rect 254791 2869 254839 2897
rect 254529 2835 254839 2869
rect 254529 2807 254577 2835
rect 254605 2807 254639 2835
rect 254667 2807 254701 2835
rect 254729 2807 254763 2835
rect 254791 2807 254839 2835
rect 254529 2773 254839 2807
rect 254529 2745 254577 2773
rect 254605 2745 254639 2773
rect 254667 2745 254701 2773
rect 254729 2745 254763 2773
rect 254791 2745 254839 2773
rect 254529 904 254839 2745
rect 254529 876 254577 904
rect 254605 876 254639 904
rect 254667 876 254701 904
rect 254729 876 254763 904
rect 254791 876 254839 904
rect 254529 842 254839 876
rect 254529 814 254577 842
rect 254605 814 254639 842
rect 254667 814 254701 842
rect 254729 814 254763 842
rect 254791 814 254839 842
rect 254529 780 254839 814
rect 254529 752 254577 780
rect 254605 752 254639 780
rect 254667 752 254701 780
rect 254729 752 254763 780
rect 254791 752 254839 780
rect 254529 718 254839 752
rect 254529 690 254577 718
rect 254605 690 254639 718
rect 254667 690 254701 718
rect 254729 690 254763 718
rect 254791 690 254839 718
rect 254529 162 254839 690
rect 256389 5959 256699 14745
rect 256389 5931 256437 5959
rect 256465 5931 256499 5959
rect 256527 5931 256561 5959
rect 256589 5931 256623 5959
rect 256651 5931 256699 5959
rect 256389 5897 256699 5931
rect 256389 5869 256437 5897
rect 256465 5869 256499 5897
rect 256527 5869 256561 5897
rect 256589 5869 256623 5897
rect 256651 5869 256699 5897
rect 256389 5835 256699 5869
rect 256389 5807 256437 5835
rect 256465 5807 256499 5835
rect 256527 5807 256561 5835
rect 256589 5807 256623 5835
rect 256651 5807 256699 5835
rect 256389 5773 256699 5807
rect 256389 5745 256437 5773
rect 256465 5745 256499 5773
rect 256527 5745 256561 5773
rect 256589 5745 256623 5773
rect 256651 5745 256699 5773
rect 256389 424 256699 5745
rect 256389 396 256437 424
rect 256465 396 256499 424
rect 256527 396 256561 424
rect 256589 396 256623 424
rect 256651 396 256699 424
rect 256389 362 256699 396
rect 256389 334 256437 362
rect 256465 334 256499 362
rect 256527 334 256561 362
rect 256589 334 256623 362
rect 256651 334 256699 362
rect 256389 300 256699 334
rect 256389 272 256437 300
rect 256465 272 256499 300
rect 256527 272 256561 300
rect 256589 272 256623 300
rect 256651 272 256699 300
rect 256389 238 256699 272
rect 256389 210 256437 238
rect 256465 210 256499 238
rect 256527 210 256561 238
rect 256589 210 256623 238
rect 256651 210 256699 238
rect 256389 162 256699 210
rect 263529 299190 263839 299718
rect 263529 299162 263577 299190
rect 263605 299162 263639 299190
rect 263667 299162 263701 299190
rect 263729 299162 263763 299190
rect 263791 299162 263839 299190
rect 263529 299128 263839 299162
rect 263529 299100 263577 299128
rect 263605 299100 263639 299128
rect 263667 299100 263701 299128
rect 263729 299100 263763 299128
rect 263791 299100 263839 299128
rect 263529 299066 263839 299100
rect 263529 299038 263577 299066
rect 263605 299038 263639 299066
rect 263667 299038 263701 299066
rect 263729 299038 263763 299066
rect 263791 299038 263839 299066
rect 263529 299004 263839 299038
rect 263529 298976 263577 299004
rect 263605 298976 263639 299004
rect 263667 298976 263701 299004
rect 263729 298976 263763 299004
rect 263791 298976 263839 299004
rect 263529 290959 263839 298976
rect 263529 290931 263577 290959
rect 263605 290931 263639 290959
rect 263667 290931 263701 290959
rect 263729 290931 263763 290959
rect 263791 290931 263839 290959
rect 263529 290897 263839 290931
rect 263529 290869 263577 290897
rect 263605 290869 263639 290897
rect 263667 290869 263701 290897
rect 263729 290869 263763 290897
rect 263791 290869 263839 290897
rect 263529 290835 263839 290869
rect 263529 290807 263577 290835
rect 263605 290807 263639 290835
rect 263667 290807 263701 290835
rect 263729 290807 263763 290835
rect 263791 290807 263839 290835
rect 263529 290773 263839 290807
rect 263529 290745 263577 290773
rect 263605 290745 263639 290773
rect 263667 290745 263701 290773
rect 263729 290745 263763 290773
rect 263791 290745 263839 290773
rect 263529 281959 263839 290745
rect 263529 281931 263577 281959
rect 263605 281931 263639 281959
rect 263667 281931 263701 281959
rect 263729 281931 263763 281959
rect 263791 281931 263839 281959
rect 263529 281897 263839 281931
rect 263529 281869 263577 281897
rect 263605 281869 263639 281897
rect 263667 281869 263701 281897
rect 263729 281869 263763 281897
rect 263791 281869 263839 281897
rect 263529 281835 263839 281869
rect 263529 281807 263577 281835
rect 263605 281807 263639 281835
rect 263667 281807 263701 281835
rect 263729 281807 263763 281835
rect 263791 281807 263839 281835
rect 263529 281773 263839 281807
rect 263529 281745 263577 281773
rect 263605 281745 263639 281773
rect 263667 281745 263701 281773
rect 263729 281745 263763 281773
rect 263791 281745 263839 281773
rect 263529 272959 263839 281745
rect 263529 272931 263577 272959
rect 263605 272931 263639 272959
rect 263667 272931 263701 272959
rect 263729 272931 263763 272959
rect 263791 272931 263839 272959
rect 263529 272897 263839 272931
rect 263529 272869 263577 272897
rect 263605 272869 263639 272897
rect 263667 272869 263701 272897
rect 263729 272869 263763 272897
rect 263791 272869 263839 272897
rect 263529 272835 263839 272869
rect 263529 272807 263577 272835
rect 263605 272807 263639 272835
rect 263667 272807 263701 272835
rect 263729 272807 263763 272835
rect 263791 272807 263839 272835
rect 263529 272773 263839 272807
rect 263529 272745 263577 272773
rect 263605 272745 263639 272773
rect 263667 272745 263701 272773
rect 263729 272745 263763 272773
rect 263791 272745 263839 272773
rect 263529 263959 263839 272745
rect 263529 263931 263577 263959
rect 263605 263931 263639 263959
rect 263667 263931 263701 263959
rect 263729 263931 263763 263959
rect 263791 263931 263839 263959
rect 263529 263897 263839 263931
rect 263529 263869 263577 263897
rect 263605 263869 263639 263897
rect 263667 263869 263701 263897
rect 263729 263869 263763 263897
rect 263791 263869 263839 263897
rect 263529 263835 263839 263869
rect 263529 263807 263577 263835
rect 263605 263807 263639 263835
rect 263667 263807 263701 263835
rect 263729 263807 263763 263835
rect 263791 263807 263839 263835
rect 263529 263773 263839 263807
rect 263529 263745 263577 263773
rect 263605 263745 263639 263773
rect 263667 263745 263701 263773
rect 263729 263745 263763 263773
rect 263791 263745 263839 263773
rect 263529 254959 263839 263745
rect 263529 254931 263577 254959
rect 263605 254931 263639 254959
rect 263667 254931 263701 254959
rect 263729 254931 263763 254959
rect 263791 254931 263839 254959
rect 263529 254897 263839 254931
rect 263529 254869 263577 254897
rect 263605 254869 263639 254897
rect 263667 254869 263701 254897
rect 263729 254869 263763 254897
rect 263791 254869 263839 254897
rect 263529 254835 263839 254869
rect 263529 254807 263577 254835
rect 263605 254807 263639 254835
rect 263667 254807 263701 254835
rect 263729 254807 263763 254835
rect 263791 254807 263839 254835
rect 263529 254773 263839 254807
rect 263529 254745 263577 254773
rect 263605 254745 263639 254773
rect 263667 254745 263701 254773
rect 263729 254745 263763 254773
rect 263791 254745 263839 254773
rect 263529 245959 263839 254745
rect 263529 245931 263577 245959
rect 263605 245931 263639 245959
rect 263667 245931 263701 245959
rect 263729 245931 263763 245959
rect 263791 245931 263839 245959
rect 263529 245897 263839 245931
rect 263529 245869 263577 245897
rect 263605 245869 263639 245897
rect 263667 245869 263701 245897
rect 263729 245869 263763 245897
rect 263791 245869 263839 245897
rect 263529 245835 263839 245869
rect 263529 245807 263577 245835
rect 263605 245807 263639 245835
rect 263667 245807 263701 245835
rect 263729 245807 263763 245835
rect 263791 245807 263839 245835
rect 263529 245773 263839 245807
rect 263529 245745 263577 245773
rect 263605 245745 263639 245773
rect 263667 245745 263701 245773
rect 263729 245745 263763 245773
rect 263791 245745 263839 245773
rect 263529 236959 263839 245745
rect 263529 236931 263577 236959
rect 263605 236931 263639 236959
rect 263667 236931 263701 236959
rect 263729 236931 263763 236959
rect 263791 236931 263839 236959
rect 263529 236897 263839 236931
rect 263529 236869 263577 236897
rect 263605 236869 263639 236897
rect 263667 236869 263701 236897
rect 263729 236869 263763 236897
rect 263791 236869 263839 236897
rect 263529 236835 263839 236869
rect 263529 236807 263577 236835
rect 263605 236807 263639 236835
rect 263667 236807 263701 236835
rect 263729 236807 263763 236835
rect 263791 236807 263839 236835
rect 263529 236773 263839 236807
rect 263529 236745 263577 236773
rect 263605 236745 263639 236773
rect 263667 236745 263701 236773
rect 263729 236745 263763 236773
rect 263791 236745 263839 236773
rect 263529 227959 263839 236745
rect 263529 227931 263577 227959
rect 263605 227931 263639 227959
rect 263667 227931 263701 227959
rect 263729 227931 263763 227959
rect 263791 227931 263839 227959
rect 263529 227897 263839 227931
rect 263529 227869 263577 227897
rect 263605 227869 263639 227897
rect 263667 227869 263701 227897
rect 263729 227869 263763 227897
rect 263791 227869 263839 227897
rect 263529 227835 263839 227869
rect 263529 227807 263577 227835
rect 263605 227807 263639 227835
rect 263667 227807 263701 227835
rect 263729 227807 263763 227835
rect 263791 227807 263839 227835
rect 263529 227773 263839 227807
rect 263529 227745 263577 227773
rect 263605 227745 263639 227773
rect 263667 227745 263701 227773
rect 263729 227745 263763 227773
rect 263791 227745 263839 227773
rect 263529 218959 263839 227745
rect 263529 218931 263577 218959
rect 263605 218931 263639 218959
rect 263667 218931 263701 218959
rect 263729 218931 263763 218959
rect 263791 218931 263839 218959
rect 263529 218897 263839 218931
rect 263529 218869 263577 218897
rect 263605 218869 263639 218897
rect 263667 218869 263701 218897
rect 263729 218869 263763 218897
rect 263791 218869 263839 218897
rect 263529 218835 263839 218869
rect 263529 218807 263577 218835
rect 263605 218807 263639 218835
rect 263667 218807 263701 218835
rect 263729 218807 263763 218835
rect 263791 218807 263839 218835
rect 263529 218773 263839 218807
rect 263529 218745 263577 218773
rect 263605 218745 263639 218773
rect 263667 218745 263701 218773
rect 263729 218745 263763 218773
rect 263791 218745 263839 218773
rect 263529 209959 263839 218745
rect 263529 209931 263577 209959
rect 263605 209931 263639 209959
rect 263667 209931 263701 209959
rect 263729 209931 263763 209959
rect 263791 209931 263839 209959
rect 263529 209897 263839 209931
rect 263529 209869 263577 209897
rect 263605 209869 263639 209897
rect 263667 209869 263701 209897
rect 263729 209869 263763 209897
rect 263791 209869 263839 209897
rect 263529 209835 263839 209869
rect 263529 209807 263577 209835
rect 263605 209807 263639 209835
rect 263667 209807 263701 209835
rect 263729 209807 263763 209835
rect 263791 209807 263839 209835
rect 263529 209773 263839 209807
rect 263529 209745 263577 209773
rect 263605 209745 263639 209773
rect 263667 209745 263701 209773
rect 263729 209745 263763 209773
rect 263791 209745 263839 209773
rect 263529 200959 263839 209745
rect 263529 200931 263577 200959
rect 263605 200931 263639 200959
rect 263667 200931 263701 200959
rect 263729 200931 263763 200959
rect 263791 200931 263839 200959
rect 263529 200897 263839 200931
rect 263529 200869 263577 200897
rect 263605 200869 263639 200897
rect 263667 200869 263701 200897
rect 263729 200869 263763 200897
rect 263791 200869 263839 200897
rect 263529 200835 263839 200869
rect 263529 200807 263577 200835
rect 263605 200807 263639 200835
rect 263667 200807 263701 200835
rect 263729 200807 263763 200835
rect 263791 200807 263839 200835
rect 263529 200773 263839 200807
rect 263529 200745 263577 200773
rect 263605 200745 263639 200773
rect 263667 200745 263701 200773
rect 263729 200745 263763 200773
rect 263791 200745 263839 200773
rect 263529 191959 263839 200745
rect 263529 191931 263577 191959
rect 263605 191931 263639 191959
rect 263667 191931 263701 191959
rect 263729 191931 263763 191959
rect 263791 191931 263839 191959
rect 263529 191897 263839 191931
rect 263529 191869 263577 191897
rect 263605 191869 263639 191897
rect 263667 191869 263701 191897
rect 263729 191869 263763 191897
rect 263791 191869 263839 191897
rect 263529 191835 263839 191869
rect 263529 191807 263577 191835
rect 263605 191807 263639 191835
rect 263667 191807 263701 191835
rect 263729 191807 263763 191835
rect 263791 191807 263839 191835
rect 263529 191773 263839 191807
rect 263529 191745 263577 191773
rect 263605 191745 263639 191773
rect 263667 191745 263701 191773
rect 263729 191745 263763 191773
rect 263791 191745 263839 191773
rect 263529 182959 263839 191745
rect 263529 182931 263577 182959
rect 263605 182931 263639 182959
rect 263667 182931 263701 182959
rect 263729 182931 263763 182959
rect 263791 182931 263839 182959
rect 263529 182897 263839 182931
rect 263529 182869 263577 182897
rect 263605 182869 263639 182897
rect 263667 182869 263701 182897
rect 263729 182869 263763 182897
rect 263791 182869 263839 182897
rect 263529 182835 263839 182869
rect 263529 182807 263577 182835
rect 263605 182807 263639 182835
rect 263667 182807 263701 182835
rect 263729 182807 263763 182835
rect 263791 182807 263839 182835
rect 263529 182773 263839 182807
rect 263529 182745 263577 182773
rect 263605 182745 263639 182773
rect 263667 182745 263701 182773
rect 263729 182745 263763 182773
rect 263791 182745 263839 182773
rect 263529 173959 263839 182745
rect 263529 173931 263577 173959
rect 263605 173931 263639 173959
rect 263667 173931 263701 173959
rect 263729 173931 263763 173959
rect 263791 173931 263839 173959
rect 263529 173897 263839 173931
rect 263529 173869 263577 173897
rect 263605 173869 263639 173897
rect 263667 173869 263701 173897
rect 263729 173869 263763 173897
rect 263791 173869 263839 173897
rect 263529 173835 263839 173869
rect 263529 173807 263577 173835
rect 263605 173807 263639 173835
rect 263667 173807 263701 173835
rect 263729 173807 263763 173835
rect 263791 173807 263839 173835
rect 263529 173773 263839 173807
rect 263529 173745 263577 173773
rect 263605 173745 263639 173773
rect 263667 173745 263701 173773
rect 263729 173745 263763 173773
rect 263791 173745 263839 173773
rect 263529 164959 263839 173745
rect 263529 164931 263577 164959
rect 263605 164931 263639 164959
rect 263667 164931 263701 164959
rect 263729 164931 263763 164959
rect 263791 164931 263839 164959
rect 263529 164897 263839 164931
rect 263529 164869 263577 164897
rect 263605 164869 263639 164897
rect 263667 164869 263701 164897
rect 263729 164869 263763 164897
rect 263791 164869 263839 164897
rect 263529 164835 263839 164869
rect 263529 164807 263577 164835
rect 263605 164807 263639 164835
rect 263667 164807 263701 164835
rect 263729 164807 263763 164835
rect 263791 164807 263839 164835
rect 263529 164773 263839 164807
rect 263529 164745 263577 164773
rect 263605 164745 263639 164773
rect 263667 164745 263701 164773
rect 263729 164745 263763 164773
rect 263791 164745 263839 164773
rect 263529 155959 263839 164745
rect 263529 155931 263577 155959
rect 263605 155931 263639 155959
rect 263667 155931 263701 155959
rect 263729 155931 263763 155959
rect 263791 155931 263839 155959
rect 263529 155897 263839 155931
rect 263529 155869 263577 155897
rect 263605 155869 263639 155897
rect 263667 155869 263701 155897
rect 263729 155869 263763 155897
rect 263791 155869 263839 155897
rect 263529 155835 263839 155869
rect 263529 155807 263577 155835
rect 263605 155807 263639 155835
rect 263667 155807 263701 155835
rect 263729 155807 263763 155835
rect 263791 155807 263839 155835
rect 263529 155773 263839 155807
rect 263529 155745 263577 155773
rect 263605 155745 263639 155773
rect 263667 155745 263701 155773
rect 263729 155745 263763 155773
rect 263791 155745 263839 155773
rect 263529 146959 263839 155745
rect 263529 146931 263577 146959
rect 263605 146931 263639 146959
rect 263667 146931 263701 146959
rect 263729 146931 263763 146959
rect 263791 146931 263839 146959
rect 263529 146897 263839 146931
rect 263529 146869 263577 146897
rect 263605 146869 263639 146897
rect 263667 146869 263701 146897
rect 263729 146869 263763 146897
rect 263791 146869 263839 146897
rect 263529 146835 263839 146869
rect 263529 146807 263577 146835
rect 263605 146807 263639 146835
rect 263667 146807 263701 146835
rect 263729 146807 263763 146835
rect 263791 146807 263839 146835
rect 263529 146773 263839 146807
rect 263529 146745 263577 146773
rect 263605 146745 263639 146773
rect 263667 146745 263701 146773
rect 263729 146745 263763 146773
rect 263791 146745 263839 146773
rect 263529 137959 263839 146745
rect 263529 137931 263577 137959
rect 263605 137931 263639 137959
rect 263667 137931 263701 137959
rect 263729 137931 263763 137959
rect 263791 137931 263839 137959
rect 263529 137897 263839 137931
rect 263529 137869 263577 137897
rect 263605 137869 263639 137897
rect 263667 137869 263701 137897
rect 263729 137869 263763 137897
rect 263791 137869 263839 137897
rect 263529 137835 263839 137869
rect 263529 137807 263577 137835
rect 263605 137807 263639 137835
rect 263667 137807 263701 137835
rect 263729 137807 263763 137835
rect 263791 137807 263839 137835
rect 263529 137773 263839 137807
rect 263529 137745 263577 137773
rect 263605 137745 263639 137773
rect 263667 137745 263701 137773
rect 263729 137745 263763 137773
rect 263791 137745 263839 137773
rect 263529 128959 263839 137745
rect 263529 128931 263577 128959
rect 263605 128931 263639 128959
rect 263667 128931 263701 128959
rect 263729 128931 263763 128959
rect 263791 128931 263839 128959
rect 263529 128897 263839 128931
rect 263529 128869 263577 128897
rect 263605 128869 263639 128897
rect 263667 128869 263701 128897
rect 263729 128869 263763 128897
rect 263791 128869 263839 128897
rect 263529 128835 263839 128869
rect 263529 128807 263577 128835
rect 263605 128807 263639 128835
rect 263667 128807 263701 128835
rect 263729 128807 263763 128835
rect 263791 128807 263839 128835
rect 263529 128773 263839 128807
rect 263529 128745 263577 128773
rect 263605 128745 263639 128773
rect 263667 128745 263701 128773
rect 263729 128745 263763 128773
rect 263791 128745 263839 128773
rect 263529 119959 263839 128745
rect 263529 119931 263577 119959
rect 263605 119931 263639 119959
rect 263667 119931 263701 119959
rect 263729 119931 263763 119959
rect 263791 119931 263839 119959
rect 263529 119897 263839 119931
rect 263529 119869 263577 119897
rect 263605 119869 263639 119897
rect 263667 119869 263701 119897
rect 263729 119869 263763 119897
rect 263791 119869 263839 119897
rect 263529 119835 263839 119869
rect 263529 119807 263577 119835
rect 263605 119807 263639 119835
rect 263667 119807 263701 119835
rect 263729 119807 263763 119835
rect 263791 119807 263839 119835
rect 263529 119773 263839 119807
rect 263529 119745 263577 119773
rect 263605 119745 263639 119773
rect 263667 119745 263701 119773
rect 263729 119745 263763 119773
rect 263791 119745 263839 119773
rect 263529 110959 263839 119745
rect 263529 110931 263577 110959
rect 263605 110931 263639 110959
rect 263667 110931 263701 110959
rect 263729 110931 263763 110959
rect 263791 110931 263839 110959
rect 263529 110897 263839 110931
rect 263529 110869 263577 110897
rect 263605 110869 263639 110897
rect 263667 110869 263701 110897
rect 263729 110869 263763 110897
rect 263791 110869 263839 110897
rect 263529 110835 263839 110869
rect 263529 110807 263577 110835
rect 263605 110807 263639 110835
rect 263667 110807 263701 110835
rect 263729 110807 263763 110835
rect 263791 110807 263839 110835
rect 263529 110773 263839 110807
rect 263529 110745 263577 110773
rect 263605 110745 263639 110773
rect 263667 110745 263701 110773
rect 263729 110745 263763 110773
rect 263791 110745 263839 110773
rect 263529 101959 263839 110745
rect 263529 101931 263577 101959
rect 263605 101931 263639 101959
rect 263667 101931 263701 101959
rect 263729 101931 263763 101959
rect 263791 101931 263839 101959
rect 263529 101897 263839 101931
rect 263529 101869 263577 101897
rect 263605 101869 263639 101897
rect 263667 101869 263701 101897
rect 263729 101869 263763 101897
rect 263791 101869 263839 101897
rect 263529 101835 263839 101869
rect 263529 101807 263577 101835
rect 263605 101807 263639 101835
rect 263667 101807 263701 101835
rect 263729 101807 263763 101835
rect 263791 101807 263839 101835
rect 263529 101773 263839 101807
rect 263529 101745 263577 101773
rect 263605 101745 263639 101773
rect 263667 101745 263701 101773
rect 263729 101745 263763 101773
rect 263791 101745 263839 101773
rect 263529 92959 263839 101745
rect 263529 92931 263577 92959
rect 263605 92931 263639 92959
rect 263667 92931 263701 92959
rect 263729 92931 263763 92959
rect 263791 92931 263839 92959
rect 263529 92897 263839 92931
rect 263529 92869 263577 92897
rect 263605 92869 263639 92897
rect 263667 92869 263701 92897
rect 263729 92869 263763 92897
rect 263791 92869 263839 92897
rect 263529 92835 263839 92869
rect 263529 92807 263577 92835
rect 263605 92807 263639 92835
rect 263667 92807 263701 92835
rect 263729 92807 263763 92835
rect 263791 92807 263839 92835
rect 263529 92773 263839 92807
rect 263529 92745 263577 92773
rect 263605 92745 263639 92773
rect 263667 92745 263701 92773
rect 263729 92745 263763 92773
rect 263791 92745 263839 92773
rect 263529 83959 263839 92745
rect 263529 83931 263577 83959
rect 263605 83931 263639 83959
rect 263667 83931 263701 83959
rect 263729 83931 263763 83959
rect 263791 83931 263839 83959
rect 263529 83897 263839 83931
rect 263529 83869 263577 83897
rect 263605 83869 263639 83897
rect 263667 83869 263701 83897
rect 263729 83869 263763 83897
rect 263791 83869 263839 83897
rect 263529 83835 263839 83869
rect 263529 83807 263577 83835
rect 263605 83807 263639 83835
rect 263667 83807 263701 83835
rect 263729 83807 263763 83835
rect 263791 83807 263839 83835
rect 263529 83773 263839 83807
rect 263529 83745 263577 83773
rect 263605 83745 263639 83773
rect 263667 83745 263701 83773
rect 263729 83745 263763 83773
rect 263791 83745 263839 83773
rect 263529 74959 263839 83745
rect 263529 74931 263577 74959
rect 263605 74931 263639 74959
rect 263667 74931 263701 74959
rect 263729 74931 263763 74959
rect 263791 74931 263839 74959
rect 263529 74897 263839 74931
rect 263529 74869 263577 74897
rect 263605 74869 263639 74897
rect 263667 74869 263701 74897
rect 263729 74869 263763 74897
rect 263791 74869 263839 74897
rect 263529 74835 263839 74869
rect 263529 74807 263577 74835
rect 263605 74807 263639 74835
rect 263667 74807 263701 74835
rect 263729 74807 263763 74835
rect 263791 74807 263839 74835
rect 263529 74773 263839 74807
rect 263529 74745 263577 74773
rect 263605 74745 263639 74773
rect 263667 74745 263701 74773
rect 263729 74745 263763 74773
rect 263791 74745 263839 74773
rect 263529 65959 263839 74745
rect 263529 65931 263577 65959
rect 263605 65931 263639 65959
rect 263667 65931 263701 65959
rect 263729 65931 263763 65959
rect 263791 65931 263839 65959
rect 263529 65897 263839 65931
rect 263529 65869 263577 65897
rect 263605 65869 263639 65897
rect 263667 65869 263701 65897
rect 263729 65869 263763 65897
rect 263791 65869 263839 65897
rect 263529 65835 263839 65869
rect 263529 65807 263577 65835
rect 263605 65807 263639 65835
rect 263667 65807 263701 65835
rect 263729 65807 263763 65835
rect 263791 65807 263839 65835
rect 263529 65773 263839 65807
rect 263529 65745 263577 65773
rect 263605 65745 263639 65773
rect 263667 65745 263701 65773
rect 263729 65745 263763 65773
rect 263791 65745 263839 65773
rect 263529 56959 263839 65745
rect 263529 56931 263577 56959
rect 263605 56931 263639 56959
rect 263667 56931 263701 56959
rect 263729 56931 263763 56959
rect 263791 56931 263839 56959
rect 263529 56897 263839 56931
rect 263529 56869 263577 56897
rect 263605 56869 263639 56897
rect 263667 56869 263701 56897
rect 263729 56869 263763 56897
rect 263791 56869 263839 56897
rect 263529 56835 263839 56869
rect 263529 56807 263577 56835
rect 263605 56807 263639 56835
rect 263667 56807 263701 56835
rect 263729 56807 263763 56835
rect 263791 56807 263839 56835
rect 263529 56773 263839 56807
rect 263529 56745 263577 56773
rect 263605 56745 263639 56773
rect 263667 56745 263701 56773
rect 263729 56745 263763 56773
rect 263791 56745 263839 56773
rect 263529 47959 263839 56745
rect 263529 47931 263577 47959
rect 263605 47931 263639 47959
rect 263667 47931 263701 47959
rect 263729 47931 263763 47959
rect 263791 47931 263839 47959
rect 263529 47897 263839 47931
rect 263529 47869 263577 47897
rect 263605 47869 263639 47897
rect 263667 47869 263701 47897
rect 263729 47869 263763 47897
rect 263791 47869 263839 47897
rect 263529 47835 263839 47869
rect 263529 47807 263577 47835
rect 263605 47807 263639 47835
rect 263667 47807 263701 47835
rect 263729 47807 263763 47835
rect 263791 47807 263839 47835
rect 263529 47773 263839 47807
rect 263529 47745 263577 47773
rect 263605 47745 263639 47773
rect 263667 47745 263701 47773
rect 263729 47745 263763 47773
rect 263791 47745 263839 47773
rect 263529 38959 263839 47745
rect 263529 38931 263577 38959
rect 263605 38931 263639 38959
rect 263667 38931 263701 38959
rect 263729 38931 263763 38959
rect 263791 38931 263839 38959
rect 263529 38897 263839 38931
rect 263529 38869 263577 38897
rect 263605 38869 263639 38897
rect 263667 38869 263701 38897
rect 263729 38869 263763 38897
rect 263791 38869 263839 38897
rect 263529 38835 263839 38869
rect 263529 38807 263577 38835
rect 263605 38807 263639 38835
rect 263667 38807 263701 38835
rect 263729 38807 263763 38835
rect 263791 38807 263839 38835
rect 263529 38773 263839 38807
rect 263529 38745 263577 38773
rect 263605 38745 263639 38773
rect 263667 38745 263701 38773
rect 263729 38745 263763 38773
rect 263791 38745 263839 38773
rect 263529 29959 263839 38745
rect 263529 29931 263577 29959
rect 263605 29931 263639 29959
rect 263667 29931 263701 29959
rect 263729 29931 263763 29959
rect 263791 29931 263839 29959
rect 263529 29897 263839 29931
rect 263529 29869 263577 29897
rect 263605 29869 263639 29897
rect 263667 29869 263701 29897
rect 263729 29869 263763 29897
rect 263791 29869 263839 29897
rect 263529 29835 263839 29869
rect 263529 29807 263577 29835
rect 263605 29807 263639 29835
rect 263667 29807 263701 29835
rect 263729 29807 263763 29835
rect 263791 29807 263839 29835
rect 263529 29773 263839 29807
rect 263529 29745 263577 29773
rect 263605 29745 263639 29773
rect 263667 29745 263701 29773
rect 263729 29745 263763 29773
rect 263791 29745 263839 29773
rect 263529 20959 263839 29745
rect 263529 20931 263577 20959
rect 263605 20931 263639 20959
rect 263667 20931 263701 20959
rect 263729 20931 263763 20959
rect 263791 20931 263839 20959
rect 263529 20897 263839 20931
rect 263529 20869 263577 20897
rect 263605 20869 263639 20897
rect 263667 20869 263701 20897
rect 263729 20869 263763 20897
rect 263791 20869 263839 20897
rect 263529 20835 263839 20869
rect 263529 20807 263577 20835
rect 263605 20807 263639 20835
rect 263667 20807 263701 20835
rect 263729 20807 263763 20835
rect 263791 20807 263839 20835
rect 263529 20773 263839 20807
rect 263529 20745 263577 20773
rect 263605 20745 263639 20773
rect 263667 20745 263701 20773
rect 263729 20745 263763 20773
rect 263791 20745 263839 20773
rect 263529 11959 263839 20745
rect 263529 11931 263577 11959
rect 263605 11931 263639 11959
rect 263667 11931 263701 11959
rect 263729 11931 263763 11959
rect 263791 11931 263839 11959
rect 263529 11897 263839 11931
rect 263529 11869 263577 11897
rect 263605 11869 263639 11897
rect 263667 11869 263701 11897
rect 263729 11869 263763 11897
rect 263791 11869 263839 11897
rect 263529 11835 263839 11869
rect 263529 11807 263577 11835
rect 263605 11807 263639 11835
rect 263667 11807 263701 11835
rect 263729 11807 263763 11835
rect 263791 11807 263839 11835
rect 263529 11773 263839 11807
rect 263529 11745 263577 11773
rect 263605 11745 263639 11773
rect 263667 11745 263701 11773
rect 263729 11745 263763 11773
rect 263791 11745 263839 11773
rect 263529 2959 263839 11745
rect 263529 2931 263577 2959
rect 263605 2931 263639 2959
rect 263667 2931 263701 2959
rect 263729 2931 263763 2959
rect 263791 2931 263839 2959
rect 263529 2897 263839 2931
rect 263529 2869 263577 2897
rect 263605 2869 263639 2897
rect 263667 2869 263701 2897
rect 263729 2869 263763 2897
rect 263791 2869 263839 2897
rect 263529 2835 263839 2869
rect 263529 2807 263577 2835
rect 263605 2807 263639 2835
rect 263667 2807 263701 2835
rect 263729 2807 263763 2835
rect 263791 2807 263839 2835
rect 263529 2773 263839 2807
rect 263529 2745 263577 2773
rect 263605 2745 263639 2773
rect 263667 2745 263701 2773
rect 263729 2745 263763 2773
rect 263791 2745 263839 2773
rect 263529 904 263839 2745
rect 263529 876 263577 904
rect 263605 876 263639 904
rect 263667 876 263701 904
rect 263729 876 263763 904
rect 263791 876 263839 904
rect 263529 842 263839 876
rect 263529 814 263577 842
rect 263605 814 263639 842
rect 263667 814 263701 842
rect 263729 814 263763 842
rect 263791 814 263839 842
rect 263529 780 263839 814
rect 263529 752 263577 780
rect 263605 752 263639 780
rect 263667 752 263701 780
rect 263729 752 263763 780
rect 263791 752 263839 780
rect 263529 718 263839 752
rect 263529 690 263577 718
rect 263605 690 263639 718
rect 263667 690 263701 718
rect 263729 690 263763 718
rect 263791 690 263839 718
rect 263529 162 263839 690
rect 265389 299670 265699 299718
rect 265389 299642 265437 299670
rect 265465 299642 265499 299670
rect 265527 299642 265561 299670
rect 265589 299642 265623 299670
rect 265651 299642 265699 299670
rect 265389 299608 265699 299642
rect 265389 299580 265437 299608
rect 265465 299580 265499 299608
rect 265527 299580 265561 299608
rect 265589 299580 265623 299608
rect 265651 299580 265699 299608
rect 265389 299546 265699 299580
rect 265389 299518 265437 299546
rect 265465 299518 265499 299546
rect 265527 299518 265561 299546
rect 265589 299518 265623 299546
rect 265651 299518 265699 299546
rect 265389 299484 265699 299518
rect 265389 299456 265437 299484
rect 265465 299456 265499 299484
rect 265527 299456 265561 299484
rect 265589 299456 265623 299484
rect 265651 299456 265699 299484
rect 265389 293959 265699 299456
rect 265389 293931 265437 293959
rect 265465 293931 265499 293959
rect 265527 293931 265561 293959
rect 265589 293931 265623 293959
rect 265651 293931 265699 293959
rect 265389 293897 265699 293931
rect 265389 293869 265437 293897
rect 265465 293869 265499 293897
rect 265527 293869 265561 293897
rect 265589 293869 265623 293897
rect 265651 293869 265699 293897
rect 265389 293835 265699 293869
rect 265389 293807 265437 293835
rect 265465 293807 265499 293835
rect 265527 293807 265561 293835
rect 265589 293807 265623 293835
rect 265651 293807 265699 293835
rect 265389 293773 265699 293807
rect 265389 293745 265437 293773
rect 265465 293745 265499 293773
rect 265527 293745 265561 293773
rect 265589 293745 265623 293773
rect 265651 293745 265699 293773
rect 265389 284959 265699 293745
rect 265389 284931 265437 284959
rect 265465 284931 265499 284959
rect 265527 284931 265561 284959
rect 265589 284931 265623 284959
rect 265651 284931 265699 284959
rect 265389 284897 265699 284931
rect 265389 284869 265437 284897
rect 265465 284869 265499 284897
rect 265527 284869 265561 284897
rect 265589 284869 265623 284897
rect 265651 284869 265699 284897
rect 265389 284835 265699 284869
rect 265389 284807 265437 284835
rect 265465 284807 265499 284835
rect 265527 284807 265561 284835
rect 265589 284807 265623 284835
rect 265651 284807 265699 284835
rect 265389 284773 265699 284807
rect 265389 284745 265437 284773
rect 265465 284745 265499 284773
rect 265527 284745 265561 284773
rect 265589 284745 265623 284773
rect 265651 284745 265699 284773
rect 265389 275959 265699 284745
rect 265389 275931 265437 275959
rect 265465 275931 265499 275959
rect 265527 275931 265561 275959
rect 265589 275931 265623 275959
rect 265651 275931 265699 275959
rect 265389 275897 265699 275931
rect 265389 275869 265437 275897
rect 265465 275869 265499 275897
rect 265527 275869 265561 275897
rect 265589 275869 265623 275897
rect 265651 275869 265699 275897
rect 265389 275835 265699 275869
rect 265389 275807 265437 275835
rect 265465 275807 265499 275835
rect 265527 275807 265561 275835
rect 265589 275807 265623 275835
rect 265651 275807 265699 275835
rect 265389 275773 265699 275807
rect 265389 275745 265437 275773
rect 265465 275745 265499 275773
rect 265527 275745 265561 275773
rect 265589 275745 265623 275773
rect 265651 275745 265699 275773
rect 265389 266959 265699 275745
rect 265389 266931 265437 266959
rect 265465 266931 265499 266959
rect 265527 266931 265561 266959
rect 265589 266931 265623 266959
rect 265651 266931 265699 266959
rect 265389 266897 265699 266931
rect 265389 266869 265437 266897
rect 265465 266869 265499 266897
rect 265527 266869 265561 266897
rect 265589 266869 265623 266897
rect 265651 266869 265699 266897
rect 265389 266835 265699 266869
rect 265389 266807 265437 266835
rect 265465 266807 265499 266835
rect 265527 266807 265561 266835
rect 265589 266807 265623 266835
rect 265651 266807 265699 266835
rect 265389 266773 265699 266807
rect 265389 266745 265437 266773
rect 265465 266745 265499 266773
rect 265527 266745 265561 266773
rect 265589 266745 265623 266773
rect 265651 266745 265699 266773
rect 265389 257959 265699 266745
rect 265389 257931 265437 257959
rect 265465 257931 265499 257959
rect 265527 257931 265561 257959
rect 265589 257931 265623 257959
rect 265651 257931 265699 257959
rect 265389 257897 265699 257931
rect 265389 257869 265437 257897
rect 265465 257869 265499 257897
rect 265527 257869 265561 257897
rect 265589 257869 265623 257897
rect 265651 257869 265699 257897
rect 265389 257835 265699 257869
rect 265389 257807 265437 257835
rect 265465 257807 265499 257835
rect 265527 257807 265561 257835
rect 265589 257807 265623 257835
rect 265651 257807 265699 257835
rect 265389 257773 265699 257807
rect 265389 257745 265437 257773
rect 265465 257745 265499 257773
rect 265527 257745 265561 257773
rect 265589 257745 265623 257773
rect 265651 257745 265699 257773
rect 265389 248959 265699 257745
rect 265389 248931 265437 248959
rect 265465 248931 265499 248959
rect 265527 248931 265561 248959
rect 265589 248931 265623 248959
rect 265651 248931 265699 248959
rect 265389 248897 265699 248931
rect 265389 248869 265437 248897
rect 265465 248869 265499 248897
rect 265527 248869 265561 248897
rect 265589 248869 265623 248897
rect 265651 248869 265699 248897
rect 265389 248835 265699 248869
rect 265389 248807 265437 248835
rect 265465 248807 265499 248835
rect 265527 248807 265561 248835
rect 265589 248807 265623 248835
rect 265651 248807 265699 248835
rect 265389 248773 265699 248807
rect 265389 248745 265437 248773
rect 265465 248745 265499 248773
rect 265527 248745 265561 248773
rect 265589 248745 265623 248773
rect 265651 248745 265699 248773
rect 265389 239959 265699 248745
rect 265389 239931 265437 239959
rect 265465 239931 265499 239959
rect 265527 239931 265561 239959
rect 265589 239931 265623 239959
rect 265651 239931 265699 239959
rect 265389 239897 265699 239931
rect 265389 239869 265437 239897
rect 265465 239869 265499 239897
rect 265527 239869 265561 239897
rect 265589 239869 265623 239897
rect 265651 239869 265699 239897
rect 265389 239835 265699 239869
rect 265389 239807 265437 239835
rect 265465 239807 265499 239835
rect 265527 239807 265561 239835
rect 265589 239807 265623 239835
rect 265651 239807 265699 239835
rect 265389 239773 265699 239807
rect 265389 239745 265437 239773
rect 265465 239745 265499 239773
rect 265527 239745 265561 239773
rect 265589 239745 265623 239773
rect 265651 239745 265699 239773
rect 265389 230959 265699 239745
rect 265389 230931 265437 230959
rect 265465 230931 265499 230959
rect 265527 230931 265561 230959
rect 265589 230931 265623 230959
rect 265651 230931 265699 230959
rect 265389 230897 265699 230931
rect 265389 230869 265437 230897
rect 265465 230869 265499 230897
rect 265527 230869 265561 230897
rect 265589 230869 265623 230897
rect 265651 230869 265699 230897
rect 265389 230835 265699 230869
rect 265389 230807 265437 230835
rect 265465 230807 265499 230835
rect 265527 230807 265561 230835
rect 265589 230807 265623 230835
rect 265651 230807 265699 230835
rect 265389 230773 265699 230807
rect 265389 230745 265437 230773
rect 265465 230745 265499 230773
rect 265527 230745 265561 230773
rect 265589 230745 265623 230773
rect 265651 230745 265699 230773
rect 265389 221959 265699 230745
rect 265389 221931 265437 221959
rect 265465 221931 265499 221959
rect 265527 221931 265561 221959
rect 265589 221931 265623 221959
rect 265651 221931 265699 221959
rect 265389 221897 265699 221931
rect 265389 221869 265437 221897
rect 265465 221869 265499 221897
rect 265527 221869 265561 221897
rect 265589 221869 265623 221897
rect 265651 221869 265699 221897
rect 265389 221835 265699 221869
rect 265389 221807 265437 221835
rect 265465 221807 265499 221835
rect 265527 221807 265561 221835
rect 265589 221807 265623 221835
rect 265651 221807 265699 221835
rect 265389 221773 265699 221807
rect 265389 221745 265437 221773
rect 265465 221745 265499 221773
rect 265527 221745 265561 221773
rect 265589 221745 265623 221773
rect 265651 221745 265699 221773
rect 265389 212959 265699 221745
rect 265389 212931 265437 212959
rect 265465 212931 265499 212959
rect 265527 212931 265561 212959
rect 265589 212931 265623 212959
rect 265651 212931 265699 212959
rect 265389 212897 265699 212931
rect 265389 212869 265437 212897
rect 265465 212869 265499 212897
rect 265527 212869 265561 212897
rect 265589 212869 265623 212897
rect 265651 212869 265699 212897
rect 265389 212835 265699 212869
rect 265389 212807 265437 212835
rect 265465 212807 265499 212835
rect 265527 212807 265561 212835
rect 265589 212807 265623 212835
rect 265651 212807 265699 212835
rect 265389 212773 265699 212807
rect 265389 212745 265437 212773
rect 265465 212745 265499 212773
rect 265527 212745 265561 212773
rect 265589 212745 265623 212773
rect 265651 212745 265699 212773
rect 265389 203959 265699 212745
rect 265389 203931 265437 203959
rect 265465 203931 265499 203959
rect 265527 203931 265561 203959
rect 265589 203931 265623 203959
rect 265651 203931 265699 203959
rect 265389 203897 265699 203931
rect 265389 203869 265437 203897
rect 265465 203869 265499 203897
rect 265527 203869 265561 203897
rect 265589 203869 265623 203897
rect 265651 203869 265699 203897
rect 265389 203835 265699 203869
rect 265389 203807 265437 203835
rect 265465 203807 265499 203835
rect 265527 203807 265561 203835
rect 265589 203807 265623 203835
rect 265651 203807 265699 203835
rect 265389 203773 265699 203807
rect 265389 203745 265437 203773
rect 265465 203745 265499 203773
rect 265527 203745 265561 203773
rect 265589 203745 265623 203773
rect 265651 203745 265699 203773
rect 265389 194959 265699 203745
rect 265389 194931 265437 194959
rect 265465 194931 265499 194959
rect 265527 194931 265561 194959
rect 265589 194931 265623 194959
rect 265651 194931 265699 194959
rect 265389 194897 265699 194931
rect 265389 194869 265437 194897
rect 265465 194869 265499 194897
rect 265527 194869 265561 194897
rect 265589 194869 265623 194897
rect 265651 194869 265699 194897
rect 265389 194835 265699 194869
rect 265389 194807 265437 194835
rect 265465 194807 265499 194835
rect 265527 194807 265561 194835
rect 265589 194807 265623 194835
rect 265651 194807 265699 194835
rect 265389 194773 265699 194807
rect 265389 194745 265437 194773
rect 265465 194745 265499 194773
rect 265527 194745 265561 194773
rect 265589 194745 265623 194773
rect 265651 194745 265699 194773
rect 265389 185959 265699 194745
rect 265389 185931 265437 185959
rect 265465 185931 265499 185959
rect 265527 185931 265561 185959
rect 265589 185931 265623 185959
rect 265651 185931 265699 185959
rect 265389 185897 265699 185931
rect 265389 185869 265437 185897
rect 265465 185869 265499 185897
rect 265527 185869 265561 185897
rect 265589 185869 265623 185897
rect 265651 185869 265699 185897
rect 265389 185835 265699 185869
rect 265389 185807 265437 185835
rect 265465 185807 265499 185835
rect 265527 185807 265561 185835
rect 265589 185807 265623 185835
rect 265651 185807 265699 185835
rect 265389 185773 265699 185807
rect 265389 185745 265437 185773
rect 265465 185745 265499 185773
rect 265527 185745 265561 185773
rect 265589 185745 265623 185773
rect 265651 185745 265699 185773
rect 265389 176959 265699 185745
rect 265389 176931 265437 176959
rect 265465 176931 265499 176959
rect 265527 176931 265561 176959
rect 265589 176931 265623 176959
rect 265651 176931 265699 176959
rect 265389 176897 265699 176931
rect 265389 176869 265437 176897
rect 265465 176869 265499 176897
rect 265527 176869 265561 176897
rect 265589 176869 265623 176897
rect 265651 176869 265699 176897
rect 265389 176835 265699 176869
rect 265389 176807 265437 176835
rect 265465 176807 265499 176835
rect 265527 176807 265561 176835
rect 265589 176807 265623 176835
rect 265651 176807 265699 176835
rect 265389 176773 265699 176807
rect 265389 176745 265437 176773
rect 265465 176745 265499 176773
rect 265527 176745 265561 176773
rect 265589 176745 265623 176773
rect 265651 176745 265699 176773
rect 265389 167959 265699 176745
rect 265389 167931 265437 167959
rect 265465 167931 265499 167959
rect 265527 167931 265561 167959
rect 265589 167931 265623 167959
rect 265651 167931 265699 167959
rect 265389 167897 265699 167931
rect 265389 167869 265437 167897
rect 265465 167869 265499 167897
rect 265527 167869 265561 167897
rect 265589 167869 265623 167897
rect 265651 167869 265699 167897
rect 265389 167835 265699 167869
rect 265389 167807 265437 167835
rect 265465 167807 265499 167835
rect 265527 167807 265561 167835
rect 265589 167807 265623 167835
rect 265651 167807 265699 167835
rect 265389 167773 265699 167807
rect 265389 167745 265437 167773
rect 265465 167745 265499 167773
rect 265527 167745 265561 167773
rect 265589 167745 265623 167773
rect 265651 167745 265699 167773
rect 265389 158959 265699 167745
rect 265389 158931 265437 158959
rect 265465 158931 265499 158959
rect 265527 158931 265561 158959
rect 265589 158931 265623 158959
rect 265651 158931 265699 158959
rect 265389 158897 265699 158931
rect 265389 158869 265437 158897
rect 265465 158869 265499 158897
rect 265527 158869 265561 158897
rect 265589 158869 265623 158897
rect 265651 158869 265699 158897
rect 265389 158835 265699 158869
rect 265389 158807 265437 158835
rect 265465 158807 265499 158835
rect 265527 158807 265561 158835
rect 265589 158807 265623 158835
rect 265651 158807 265699 158835
rect 265389 158773 265699 158807
rect 265389 158745 265437 158773
rect 265465 158745 265499 158773
rect 265527 158745 265561 158773
rect 265589 158745 265623 158773
rect 265651 158745 265699 158773
rect 265389 149959 265699 158745
rect 265389 149931 265437 149959
rect 265465 149931 265499 149959
rect 265527 149931 265561 149959
rect 265589 149931 265623 149959
rect 265651 149931 265699 149959
rect 265389 149897 265699 149931
rect 265389 149869 265437 149897
rect 265465 149869 265499 149897
rect 265527 149869 265561 149897
rect 265589 149869 265623 149897
rect 265651 149869 265699 149897
rect 265389 149835 265699 149869
rect 265389 149807 265437 149835
rect 265465 149807 265499 149835
rect 265527 149807 265561 149835
rect 265589 149807 265623 149835
rect 265651 149807 265699 149835
rect 265389 149773 265699 149807
rect 265389 149745 265437 149773
rect 265465 149745 265499 149773
rect 265527 149745 265561 149773
rect 265589 149745 265623 149773
rect 265651 149745 265699 149773
rect 265389 140959 265699 149745
rect 265389 140931 265437 140959
rect 265465 140931 265499 140959
rect 265527 140931 265561 140959
rect 265589 140931 265623 140959
rect 265651 140931 265699 140959
rect 265389 140897 265699 140931
rect 265389 140869 265437 140897
rect 265465 140869 265499 140897
rect 265527 140869 265561 140897
rect 265589 140869 265623 140897
rect 265651 140869 265699 140897
rect 265389 140835 265699 140869
rect 265389 140807 265437 140835
rect 265465 140807 265499 140835
rect 265527 140807 265561 140835
rect 265589 140807 265623 140835
rect 265651 140807 265699 140835
rect 265389 140773 265699 140807
rect 265389 140745 265437 140773
rect 265465 140745 265499 140773
rect 265527 140745 265561 140773
rect 265589 140745 265623 140773
rect 265651 140745 265699 140773
rect 265389 131959 265699 140745
rect 265389 131931 265437 131959
rect 265465 131931 265499 131959
rect 265527 131931 265561 131959
rect 265589 131931 265623 131959
rect 265651 131931 265699 131959
rect 265389 131897 265699 131931
rect 265389 131869 265437 131897
rect 265465 131869 265499 131897
rect 265527 131869 265561 131897
rect 265589 131869 265623 131897
rect 265651 131869 265699 131897
rect 265389 131835 265699 131869
rect 265389 131807 265437 131835
rect 265465 131807 265499 131835
rect 265527 131807 265561 131835
rect 265589 131807 265623 131835
rect 265651 131807 265699 131835
rect 265389 131773 265699 131807
rect 265389 131745 265437 131773
rect 265465 131745 265499 131773
rect 265527 131745 265561 131773
rect 265589 131745 265623 131773
rect 265651 131745 265699 131773
rect 265389 122959 265699 131745
rect 265389 122931 265437 122959
rect 265465 122931 265499 122959
rect 265527 122931 265561 122959
rect 265589 122931 265623 122959
rect 265651 122931 265699 122959
rect 265389 122897 265699 122931
rect 265389 122869 265437 122897
rect 265465 122869 265499 122897
rect 265527 122869 265561 122897
rect 265589 122869 265623 122897
rect 265651 122869 265699 122897
rect 265389 122835 265699 122869
rect 265389 122807 265437 122835
rect 265465 122807 265499 122835
rect 265527 122807 265561 122835
rect 265589 122807 265623 122835
rect 265651 122807 265699 122835
rect 265389 122773 265699 122807
rect 265389 122745 265437 122773
rect 265465 122745 265499 122773
rect 265527 122745 265561 122773
rect 265589 122745 265623 122773
rect 265651 122745 265699 122773
rect 265389 113959 265699 122745
rect 265389 113931 265437 113959
rect 265465 113931 265499 113959
rect 265527 113931 265561 113959
rect 265589 113931 265623 113959
rect 265651 113931 265699 113959
rect 265389 113897 265699 113931
rect 265389 113869 265437 113897
rect 265465 113869 265499 113897
rect 265527 113869 265561 113897
rect 265589 113869 265623 113897
rect 265651 113869 265699 113897
rect 265389 113835 265699 113869
rect 265389 113807 265437 113835
rect 265465 113807 265499 113835
rect 265527 113807 265561 113835
rect 265589 113807 265623 113835
rect 265651 113807 265699 113835
rect 265389 113773 265699 113807
rect 265389 113745 265437 113773
rect 265465 113745 265499 113773
rect 265527 113745 265561 113773
rect 265589 113745 265623 113773
rect 265651 113745 265699 113773
rect 265389 104959 265699 113745
rect 265389 104931 265437 104959
rect 265465 104931 265499 104959
rect 265527 104931 265561 104959
rect 265589 104931 265623 104959
rect 265651 104931 265699 104959
rect 265389 104897 265699 104931
rect 265389 104869 265437 104897
rect 265465 104869 265499 104897
rect 265527 104869 265561 104897
rect 265589 104869 265623 104897
rect 265651 104869 265699 104897
rect 265389 104835 265699 104869
rect 265389 104807 265437 104835
rect 265465 104807 265499 104835
rect 265527 104807 265561 104835
rect 265589 104807 265623 104835
rect 265651 104807 265699 104835
rect 265389 104773 265699 104807
rect 265389 104745 265437 104773
rect 265465 104745 265499 104773
rect 265527 104745 265561 104773
rect 265589 104745 265623 104773
rect 265651 104745 265699 104773
rect 265389 95959 265699 104745
rect 265389 95931 265437 95959
rect 265465 95931 265499 95959
rect 265527 95931 265561 95959
rect 265589 95931 265623 95959
rect 265651 95931 265699 95959
rect 265389 95897 265699 95931
rect 265389 95869 265437 95897
rect 265465 95869 265499 95897
rect 265527 95869 265561 95897
rect 265589 95869 265623 95897
rect 265651 95869 265699 95897
rect 265389 95835 265699 95869
rect 265389 95807 265437 95835
rect 265465 95807 265499 95835
rect 265527 95807 265561 95835
rect 265589 95807 265623 95835
rect 265651 95807 265699 95835
rect 265389 95773 265699 95807
rect 265389 95745 265437 95773
rect 265465 95745 265499 95773
rect 265527 95745 265561 95773
rect 265589 95745 265623 95773
rect 265651 95745 265699 95773
rect 265389 86959 265699 95745
rect 265389 86931 265437 86959
rect 265465 86931 265499 86959
rect 265527 86931 265561 86959
rect 265589 86931 265623 86959
rect 265651 86931 265699 86959
rect 265389 86897 265699 86931
rect 265389 86869 265437 86897
rect 265465 86869 265499 86897
rect 265527 86869 265561 86897
rect 265589 86869 265623 86897
rect 265651 86869 265699 86897
rect 265389 86835 265699 86869
rect 265389 86807 265437 86835
rect 265465 86807 265499 86835
rect 265527 86807 265561 86835
rect 265589 86807 265623 86835
rect 265651 86807 265699 86835
rect 265389 86773 265699 86807
rect 265389 86745 265437 86773
rect 265465 86745 265499 86773
rect 265527 86745 265561 86773
rect 265589 86745 265623 86773
rect 265651 86745 265699 86773
rect 265389 77959 265699 86745
rect 265389 77931 265437 77959
rect 265465 77931 265499 77959
rect 265527 77931 265561 77959
rect 265589 77931 265623 77959
rect 265651 77931 265699 77959
rect 265389 77897 265699 77931
rect 265389 77869 265437 77897
rect 265465 77869 265499 77897
rect 265527 77869 265561 77897
rect 265589 77869 265623 77897
rect 265651 77869 265699 77897
rect 265389 77835 265699 77869
rect 265389 77807 265437 77835
rect 265465 77807 265499 77835
rect 265527 77807 265561 77835
rect 265589 77807 265623 77835
rect 265651 77807 265699 77835
rect 265389 77773 265699 77807
rect 265389 77745 265437 77773
rect 265465 77745 265499 77773
rect 265527 77745 265561 77773
rect 265589 77745 265623 77773
rect 265651 77745 265699 77773
rect 265389 68959 265699 77745
rect 265389 68931 265437 68959
rect 265465 68931 265499 68959
rect 265527 68931 265561 68959
rect 265589 68931 265623 68959
rect 265651 68931 265699 68959
rect 265389 68897 265699 68931
rect 265389 68869 265437 68897
rect 265465 68869 265499 68897
rect 265527 68869 265561 68897
rect 265589 68869 265623 68897
rect 265651 68869 265699 68897
rect 265389 68835 265699 68869
rect 265389 68807 265437 68835
rect 265465 68807 265499 68835
rect 265527 68807 265561 68835
rect 265589 68807 265623 68835
rect 265651 68807 265699 68835
rect 265389 68773 265699 68807
rect 265389 68745 265437 68773
rect 265465 68745 265499 68773
rect 265527 68745 265561 68773
rect 265589 68745 265623 68773
rect 265651 68745 265699 68773
rect 265389 59959 265699 68745
rect 265389 59931 265437 59959
rect 265465 59931 265499 59959
rect 265527 59931 265561 59959
rect 265589 59931 265623 59959
rect 265651 59931 265699 59959
rect 265389 59897 265699 59931
rect 265389 59869 265437 59897
rect 265465 59869 265499 59897
rect 265527 59869 265561 59897
rect 265589 59869 265623 59897
rect 265651 59869 265699 59897
rect 265389 59835 265699 59869
rect 265389 59807 265437 59835
rect 265465 59807 265499 59835
rect 265527 59807 265561 59835
rect 265589 59807 265623 59835
rect 265651 59807 265699 59835
rect 265389 59773 265699 59807
rect 265389 59745 265437 59773
rect 265465 59745 265499 59773
rect 265527 59745 265561 59773
rect 265589 59745 265623 59773
rect 265651 59745 265699 59773
rect 265389 50959 265699 59745
rect 265389 50931 265437 50959
rect 265465 50931 265499 50959
rect 265527 50931 265561 50959
rect 265589 50931 265623 50959
rect 265651 50931 265699 50959
rect 265389 50897 265699 50931
rect 265389 50869 265437 50897
rect 265465 50869 265499 50897
rect 265527 50869 265561 50897
rect 265589 50869 265623 50897
rect 265651 50869 265699 50897
rect 265389 50835 265699 50869
rect 265389 50807 265437 50835
rect 265465 50807 265499 50835
rect 265527 50807 265561 50835
rect 265589 50807 265623 50835
rect 265651 50807 265699 50835
rect 265389 50773 265699 50807
rect 265389 50745 265437 50773
rect 265465 50745 265499 50773
rect 265527 50745 265561 50773
rect 265589 50745 265623 50773
rect 265651 50745 265699 50773
rect 265389 41959 265699 50745
rect 265389 41931 265437 41959
rect 265465 41931 265499 41959
rect 265527 41931 265561 41959
rect 265589 41931 265623 41959
rect 265651 41931 265699 41959
rect 265389 41897 265699 41931
rect 265389 41869 265437 41897
rect 265465 41869 265499 41897
rect 265527 41869 265561 41897
rect 265589 41869 265623 41897
rect 265651 41869 265699 41897
rect 265389 41835 265699 41869
rect 265389 41807 265437 41835
rect 265465 41807 265499 41835
rect 265527 41807 265561 41835
rect 265589 41807 265623 41835
rect 265651 41807 265699 41835
rect 265389 41773 265699 41807
rect 265389 41745 265437 41773
rect 265465 41745 265499 41773
rect 265527 41745 265561 41773
rect 265589 41745 265623 41773
rect 265651 41745 265699 41773
rect 265389 32959 265699 41745
rect 265389 32931 265437 32959
rect 265465 32931 265499 32959
rect 265527 32931 265561 32959
rect 265589 32931 265623 32959
rect 265651 32931 265699 32959
rect 265389 32897 265699 32931
rect 265389 32869 265437 32897
rect 265465 32869 265499 32897
rect 265527 32869 265561 32897
rect 265589 32869 265623 32897
rect 265651 32869 265699 32897
rect 265389 32835 265699 32869
rect 265389 32807 265437 32835
rect 265465 32807 265499 32835
rect 265527 32807 265561 32835
rect 265589 32807 265623 32835
rect 265651 32807 265699 32835
rect 265389 32773 265699 32807
rect 265389 32745 265437 32773
rect 265465 32745 265499 32773
rect 265527 32745 265561 32773
rect 265589 32745 265623 32773
rect 265651 32745 265699 32773
rect 265389 23959 265699 32745
rect 265389 23931 265437 23959
rect 265465 23931 265499 23959
rect 265527 23931 265561 23959
rect 265589 23931 265623 23959
rect 265651 23931 265699 23959
rect 265389 23897 265699 23931
rect 265389 23869 265437 23897
rect 265465 23869 265499 23897
rect 265527 23869 265561 23897
rect 265589 23869 265623 23897
rect 265651 23869 265699 23897
rect 265389 23835 265699 23869
rect 265389 23807 265437 23835
rect 265465 23807 265499 23835
rect 265527 23807 265561 23835
rect 265589 23807 265623 23835
rect 265651 23807 265699 23835
rect 265389 23773 265699 23807
rect 265389 23745 265437 23773
rect 265465 23745 265499 23773
rect 265527 23745 265561 23773
rect 265589 23745 265623 23773
rect 265651 23745 265699 23773
rect 265389 14959 265699 23745
rect 265389 14931 265437 14959
rect 265465 14931 265499 14959
rect 265527 14931 265561 14959
rect 265589 14931 265623 14959
rect 265651 14931 265699 14959
rect 265389 14897 265699 14931
rect 265389 14869 265437 14897
rect 265465 14869 265499 14897
rect 265527 14869 265561 14897
rect 265589 14869 265623 14897
rect 265651 14869 265699 14897
rect 265389 14835 265699 14869
rect 265389 14807 265437 14835
rect 265465 14807 265499 14835
rect 265527 14807 265561 14835
rect 265589 14807 265623 14835
rect 265651 14807 265699 14835
rect 265389 14773 265699 14807
rect 265389 14745 265437 14773
rect 265465 14745 265499 14773
rect 265527 14745 265561 14773
rect 265589 14745 265623 14773
rect 265651 14745 265699 14773
rect 265389 5959 265699 14745
rect 265389 5931 265437 5959
rect 265465 5931 265499 5959
rect 265527 5931 265561 5959
rect 265589 5931 265623 5959
rect 265651 5931 265699 5959
rect 265389 5897 265699 5931
rect 265389 5869 265437 5897
rect 265465 5869 265499 5897
rect 265527 5869 265561 5897
rect 265589 5869 265623 5897
rect 265651 5869 265699 5897
rect 265389 5835 265699 5869
rect 265389 5807 265437 5835
rect 265465 5807 265499 5835
rect 265527 5807 265561 5835
rect 265589 5807 265623 5835
rect 265651 5807 265699 5835
rect 265389 5773 265699 5807
rect 265389 5745 265437 5773
rect 265465 5745 265499 5773
rect 265527 5745 265561 5773
rect 265589 5745 265623 5773
rect 265651 5745 265699 5773
rect 265389 424 265699 5745
rect 265389 396 265437 424
rect 265465 396 265499 424
rect 265527 396 265561 424
rect 265589 396 265623 424
rect 265651 396 265699 424
rect 265389 362 265699 396
rect 265389 334 265437 362
rect 265465 334 265499 362
rect 265527 334 265561 362
rect 265589 334 265623 362
rect 265651 334 265699 362
rect 265389 300 265699 334
rect 265389 272 265437 300
rect 265465 272 265499 300
rect 265527 272 265561 300
rect 265589 272 265623 300
rect 265651 272 265699 300
rect 265389 238 265699 272
rect 265389 210 265437 238
rect 265465 210 265499 238
rect 265527 210 265561 238
rect 265589 210 265623 238
rect 265651 210 265699 238
rect 265389 162 265699 210
rect 272529 299190 272839 299718
rect 272529 299162 272577 299190
rect 272605 299162 272639 299190
rect 272667 299162 272701 299190
rect 272729 299162 272763 299190
rect 272791 299162 272839 299190
rect 272529 299128 272839 299162
rect 272529 299100 272577 299128
rect 272605 299100 272639 299128
rect 272667 299100 272701 299128
rect 272729 299100 272763 299128
rect 272791 299100 272839 299128
rect 272529 299066 272839 299100
rect 272529 299038 272577 299066
rect 272605 299038 272639 299066
rect 272667 299038 272701 299066
rect 272729 299038 272763 299066
rect 272791 299038 272839 299066
rect 272529 299004 272839 299038
rect 272529 298976 272577 299004
rect 272605 298976 272639 299004
rect 272667 298976 272701 299004
rect 272729 298976 272763 299004
rect 272791 298976 272839 299004
rect 272529 290959 272839 298976
rect 272529 290931 272577 290959
rect 272605 290931 272639 290959
rect 272667 290931 272701 290959
rect 272729 290931 272763 290959
rect 272791 290931 272839 290959
rect 272529 290897 272839 290931
rect 272529 290869 272577 290897
rect 272605 290869 272639 290897
rect 272667 290869 272701 290897
rect 272729 290869 272763 290897
rect 272791 290869 272839 290897
rect 272529 290835 272839 290869
rect 272529 290807 272577 290835
rect 272605 290807 272639 290835
rect 272667 290807 272701 290835
rect 272729 290807 272763 290835
rect 272791 290807 272839 290835
rect 272529 290773 272839 290807
rect 272529 290745 272577 290773
rect 272605 290745 272639 290773
rect 272667 290745 272701 290773
rect 272729 290745 272763 290773
rect 272791 290745 272839 290773
rect 272529 281959 272839 290745
rect 272529 281931 272577 281959
rect 272605 281931 272639 281959
rect 272667 281931 272701 281959
rect 272729 281931 272763 281959
rect 272791 281931 272839 281959
rect 272529 281897 272839 281931
rect 272529 281869 272577 281897
rect 272605 281869 272639 281897
rect 272667 281869 272701 281897
rect 272729 281869 272763 281897
rect 272791 281869 272839 281897
rect 272529 281835 272839 281869
rect 272529 281807 272577 281835
rect 272605 281807 272639 281835
rect 272667 281807 272701 281835
rect 272729 281807 272763 281835
rect 272791 281807 272839 281835
rect 272529 281773 272839 281807
rect 272529 281745 272577 281773
rect 272605 281745 272639 281773
rect 272667 281745 272701 281773
rect 272729 281745 272763 281773
rect 272791 281745 272839 281773
rect 272529 272959 272839 281745
rect 272529 272931 272577 272959
rect 272605 272931 272639 272959
rect 272667 272931 272701 272959
rect 272729 272931 272763 272959
rect 272791 272931 272839 272959
rect 272529 272897 272839 272931
rect 272529 272869 272577 272897
rect 272605 272869 272639 272897
rect 272667 272869 272701 272897
rect 272729 272869 272763 272897
rect 272791 272869 272839 272897
rect 272529 272835 272839 272869
rect 272529 272807 272577 272835
rect 272605 272807 272639 272835
rect 272667 272807 272701 272835
rect 272729 272807 272763 272835
rect 272791 272807 272839 272835
rect 272529 272773 272839 272807
rect 272529 272745 272577 272773
rect 272605 272745 272639 272773
rect 272667 272745 272701 272773
rect 272729 272745 272763 272773
rect 272791 272745 272839 272773
rect 272529 263959 272839 272745
rect 272529 263931 272577 263959
rect 272605 263931 272639 263959
rect 272667 263931 272701 263959
rect 272729 263931 272763 263959
rect 272791 263931 272839 263959
rect 272529 263897 272839 263931
rect 272529 263869 272577 263897
rect 272605 263869 272639 263897
rect 272667 263869 272701 263897
rect 272729 263869 272763 263897
rect 272791 263869 272839 263897
rect 272529 263835 272839 263869
rect 272529 263807 272577 263835
rect 272605 263807 272639 263835
rect 272667 263807 272701 263835
rect 272729 263807 272763 263835
rect 272791 263807 272839 263835
rect 272529 263773 272839 263807
rect 272529 263745 272577 263773
rect 272605 263745 272639 263773
rect 272667 263745 272701 263773
rect 272729 263745 272763 263773
rect 272791 263745 272839 263773
rect 272529 254959 272839 263745
rect 272529 254931 272577 254959
rect 272605 254931 272639 254959
rect 272667 254931 272701 254959
rect 272729 254931 272763 254959
rect 272791 254931 272839 254959
rect 272529 254897 272839 254931
rect 272529 254869 272577 254897
rect 272605 254869 272639 254897
rect 272667 254869 272701 254897
rect 272729 254869 272763 254897
rect 272791 254869 272839 254897
rect 272529 254835 272839 254869
rect 272529 254807 272577 254835
rect 272605 254807 272639 254835
rect 272667 254807 272701 254835
rect 272729 254807 272763 254835
rect 272791 254807 272839 254835
rect 272529 254773 272839 254807
rect 272529 254745 272577 254773
rect 272605 254745 272639 254773
rect 272667 254745 272701 254773
rect 272729 254745 272763 254773
rect 272791 254745 272839 254773
rect 272529 245959 272839 254745
rect 272529 245931 272577 245959
rect 272605 245931 272639 245959
rect 272667 245931 272701 245959
rect 272729 245931 272763 245959
rect 272791 245931 272839 245959
rect 272529 245897 272839 245931
rect 272529 245869 272577 245897
rect 272605 245869 272639 245897
rect 272667 245869 272701 245897
rect 272729 245869 272763 245897
rect 272791 245869 272839 245897
rect 272529 245835 272839 245869
rect 272529 245807 272577 245835
rect 272605 245807 272639 245835
rect 272667 245807 272701 245835
rect 272729 245807 272763 245835
rect 272791 245807 272839 245835
rect 272529 245773 272839 245807
rect 272529 245745 272577 245773
rect 272605 245745 272639 245773
rect 272667 245745 272701 245773
rect 272729 245745 272763 245773
rect 272791 245745 272839 245773
rect 272529 236959 272839 245745
rect 272529 236931 272577 236959
rect 272605 236931 272639 236959
rect 272667 236931 272701 236959
rect 272729 236931 272763 236959
rect 272791 236931 272839 236959
rect 272529 236897 272839 236931
rect 272529 236869 272577 236897
rect 272605 236869 272639 236897
rect 272667 236869 272701 236897
rect 272729 236869 272763 236897
rect 272791 236869 272839 236897
rect 272529 236835 272839 236869
rect 272529 236807 272577 236835
rect 272605 236807 272639 236835
rect 272667 236807 272701 236835
rect 272729 236807 272763 236835
rect 272791 236807 272839 236835
rect 272529 236773 272839 236807
rect 272529 236745 272577 236773
rect 272605 236745 272639 236773
rect 272667 236745 272701 236773
rect 272729 236745 272763 236773
rect 272791 236745 272839 236773
rect 272529 227959 272839 236745
rect 272529 227931 272577 227959
rect 272605 227931 272639 227959
rect 272667 227931 272701 227959
rect 272729 227931 272763 227959
rect 272791 227931 272839 227959
rect 272529 227897 272839 227931
rect 272529 227869 272577 227897
rect 272605 227869 272639 227897
rect 272667 227869 272701 227897
rect 272729 227869 272763 227897
rect 272791 227869 272839 227897
rect 272529 227835 272839 227869
rect 272529 227807 272577 227835
rect 272605 227807 272639 227835
rect 272667 227807 272701 227835
rect 272729 227807 272763 227835
rect 272791 227807 272839 227835
rect 272529 227773 272839 227807
rect 272529 227745 272577 227773
rect 272605 227745 272639 227773
rect 272667 227745 272701 227773
rect 272729 227745 272763 227773
rect 272791 227745 272839 227773
rect 272529 218959 272839 227745
rect 272529 218931 272577 218959
rect 272605 218931 272639 218959
rect 272667 218931 272701 218959
rect 272729 218931 272763 218959
rect 272791 218931 272839 218959
rect 272529 218897 272839 218931
rect 272529 218869 272577 218897
rect 272605 218869 272639 218897
rect 272667 218869 272701 218897
rect 272729 218869 272763 218897
rect 272791 218869 272839 218897
rect 272529 218835 272839 218869
rect 272529 218807 272577 218835
rect 272605 218807 272639 218835
rect 272667 218807 272701 218835
rect 272729 218807 272763 218835
rect 272791 218807 272839 218835
rect 272529 218773 272839 218807
rect 272529 218745 272577 218773
rect 272605 218745 272639 218773
rect 272667 218745 272701 218773
rect 272729 218745 272763 218773
rect 272791 218745 272839 218773
rect 272529 209959 272839 218745
rect 272529 209931 272577 209959
rect 272605 209931 272639 209959
rect 272667 209931 272701 209959
rect 272729 209931 272763 209959
rect 272791 209931 272839 209959
rect 272529 209897 272839 209931
rect 272529 209869 272577 209897
rect 272605 209869 272639 209897
rect 272667 209869 272701 209897
rect 272729 209869 272763 209897
rect 272791 209869 272839 209897
rect 272529 209835 272839 209869
rect 272529 209807 272577 209835
rect 272605 209807 272639 209835
rect 272667 209807 272701 209835
rect 272729 209807 272763 209835
rect 272791 209807 272839 209835
rect 272529 209773 272839 209807
rect 272529 209745 272577 209773
rect 272605 209745 272639 209773
rect 272667 209745 272701 209773
rect 272729 209745 272763 209773
rect 272791 209745 272839 209773
rect 272529 200959 272839 209745
rect 272529 200931 272577 200959
rect 272605 200931 272639 200959
rect 272667 200931 272701 200959
rect 272729 200931 272763 200959
rect 272791 200931 272839 200959
rect 272529 200897 272839 200931
rect 272529 200869 272577 200897
rect 272605 200869 272639 200897
rect 272667 200869 272701 200897
rect 272729 200869 272763 200897
rect 272791 200869 272839 200897
rect 272529 200835 272839 200869
rect 272529 200807 272577 200835
rect 272605 200807 272639 200835
rect 272667 200807 272701 200835
rect 272729 200807 272763 200835
rect 272791 200807 272839 200835
rect 272529 200773 272839 200807
rect 272529 200745 272577 200773
rect 272605 200745 272639 200773
rect 272667 200745 272701 200773
rect 272729 200745 272763 200773
rect 272791 200745 272839 200773
rect 272529 191959 272839 200745
rect 272529 191931 272577 191959
rect 272605 191931 272639 191959
rect 272667 191931 272701 191959
rect 272729 191931 272763 191959
rect 272791 191931 272839 191959
rect 272529 191897 272839 191931
rect 272529 191869 272577 191897
rect 272605 191869 272639 191897
rect 272667 191869 272701 191897
rect 272729 191869 272763 191897
rect 272791 191869 272839 191897
rect 272529 191835 272839 191869
rect 272529 191807 272577 191835
rect 272605 191807 272639 191835
rect 272667 191807 272701 191835
rect 272729 191807 272763 191835
rect 272791 191807 272839 191835
rect 272529 191773 272839 191807
rect 272529 191745 272577 191773
rect 272605 191745 272639 191773
rect 272667 191745 272701 191773
rect 272729 191745 272763 191773
rect 272791 191745 272839 191773
rect 272529 182959 272839 191745
rect 272529 182931 272577 182959
rect 272605 182931 272639 182959
rect 272667 182931 272701 182959
rect 272729 182931 272763 182959
rect 272791 182931 272839 182959
rect 272529 182897 272839 182931
rect 272529 182869 272577 182897
rect 272605 182869 272639 182897
rect 272667 182869 272701 182897
rect 272729 182869 272763 182897
rect 272791 182869 272839 182897
rect 272529 182835 272839 182869
rect 272529 182807 272577 182835
rect 272605 182807 272639 182835
rect 272667 182807 272701 182835
rect 272729 182807 272763 182835
rect 272791 182807 272839 182835
rect 272529 182773 272839 182807
rect 272529 182745 272577 182773
rect 272605 182745 272639 182773
rect 272667 182745 272701 182773
rect 272729 182745 272763 182773
rect 272791 182745 272839 182773
rect 272529 173959 272839 182745
rect 272529 173931 272577 173959
rect 272605 173931 272639 173959
rect 272667 173931 272701 173959
rect 272729 173931 272763 173959
rect 272791 173931 272839 173959
rect 272529 173897 272839 173931
rect 272529 173869 272577 173897
rect 272605 173869 272639 173897
rect 272667 173869 272701 173897
rect 272729 173869 272763 173897
rect 272791 173869 272839 173897
rect 272529 173835 272839 173869
rect 272529 173807 272577 173835
rect 272605 173807 272639 173835
rect 272667 173807 272701 173835
rect 272729 173807 272763 173835
rect 272791 173807 272839 173835
rect 272529 173773 272839 173807
rect 272529 173745 272577 173773
rect 272605 173745 272639 173773
rect 272667 173745 272701 173773
rect 272729 173745 272763 173773
rect 272791 173745 272839 173773
rect 272529 164959 272839 173745
rect 272529 164931 272577 164959
rect 272605 164931 272639 164959
rect 272667 164931 272701 164959
rect 272729 164931 272763 164959
rect 272791 164931 272839 164959
rect 272529 164897 272839 164931
rect 272529 164869 272577 164897
rect 272605 164869 272639 164897
rect 272667 164869 272701 164897
rect 272729 164869 272763 164897
rect 272791 164869 272839 164897
rect 272529 164835 272839 164869
rect 272529 164807 272577 164835
rect 272605 164807 272639 164835
rect 272667 164807 272701 164835
rect 272729 164807 272763 164835
rect 272791 164807 272839 164835
rect 272529 164773 272839 164807
rect 272529 164745 272577 164773
rect 272605 164745 272639 164773
rect 272667 164745 272701 164773
rect 272729 164745 272763 164773
rect 272791 164745 272839 164773
rect 272529 155959 272839 164745
rect 272529 155931 272577 155959
rect 272605 155931 272639 155959
rect 272667 155931 272701 155959
rect 272729 155931 272763 155959
rect 272791 155931 272839 155959
rect 272529 155897 272839 155931
rect 272529 155869 272577 155897
rect 272605 155869 272639 155897
rect 272667 155869 272701 155897
rect 272729 155869 272763 155897
rect 272791 155869 272839 155897
rect 272529 155835 272839 155869
rect 272529 155807 272577 155835
rect 272605 155807 272639 155835
rect 272667 155807 272701 155835
rect 272729 155807 272763 155835
rect 272791 155807 272839 155835
rect 272529 155773 272839 155807
rect 272529 155745 272577 155773
rect 272605 155745 272639 155773
rect 272667 155745 272701 155773
rect 272729 155745 272763 155773
rect 272791 155745 272839 155773
rect 272529 146959 272839 155745
rect 272529 146931 272577 146959
rect 272605 146931 272639 146959
rect 272667 146931 272701 146959
rect 272729 146931 272763 146959
rect 272791 146931 272839 146959
rect 272529 146897 272839 146931
rect 272529 146869 272577 146897
rect 272605 146869 272639 146897
rect 272667 146869 272701 146897
rect 272729 146869 272763 146897
rect 272791 146869 272839 146897
rect 272529 146835 272839 146869
rect 272529 146807 272577 146835
rect 272605 146807 272639 146835
rect 272667 146807 272701 146835
rect 272729 146807 272763 146835
rect 272791 146807 272839 146835
rect 272529 146773 272839 146807
rect 272529 146745 272577 146773
rect 272605 146745 272639 146773
rect 272667 146745 272701 146773
rect 272729 146745 272763 146773
rect 272791 146745 272839 146773
rect 272529 137959 272839 146745
rect 272529 137931 272577 137959
rect 272605 137931 272639 137959
rect 272667 137931 272701 137959
rect 272729 137931 272763 137959
rect 272791 137931 272839 137959
rect 272529 137897 272839 137931
rect 272529 137869 272577 137897
rect 272605 137869 272639 137897
rect 272667 137869 272701 137897
rect 272729 137869 272763 137897
rect 272791 137869 272839 137897
rect 272529 137835 272839 137869
rect 272529 137807 272577 137835
rect 272605 137807 272639 137835
rect 272667 137807 272701 137835
rect 272729 137807 272763 137835
rect 272791 137807 272839 137835
rect 272529 137773 272839 137807
rect 272529 137745 272577 137773
rect 272605 137745 272639 137773
rect 272667 137745 272701 137773
rect 272729 137745 272763 137773
rect 272791 137745 272839 137773
rect 272529 128959 272839 137745
rect 272529 128931 272577 128959
rect 272605 128931 272639 128959
rect 272667 128931 272701 128959
rect 272729 128931 272763 128959
rect 272791 128931 272839 128959
rect 272529 128897 272839 128931
rect 272529 128869 272577 128897
rect 272605 128869 272639 128897
rect 272667 128869 272701 128897
rect 272729 128869 272763 128897
rect 272791 128869 272839 128897
rect 272529 128835 272839 128869
rect 272529 128807 272577 128835
rect 272605 128807 272639 128835
rect 272667 128807 272701 128835
rect 272729 128807 272763 128835
rect 272791 128807 272839 128835
rect 272529 128773 272839 128807
rect 272529 128745 272577 128773
rect 272605 128745 272639 128773
rect 272667 128745 272701 128773
rect 272729 128745 272763 128773
rect 272791 128745 272839 128773
rect 272529 119959 272839 128745
rect 272529 119931 272577 119959
rect 272605 119931 272639 119959
rect 272667 119931 272701 119959
rect 272729 119931 272763 119959
rect 272791 119931 272839 119959
rect 272529 119897 272839 119931
rect 272529 119869 272577 119897
rect 272605 119869 272639 119897
rect 272667 119869 272701 119897
rect 272729 119869 272763 119897
rect 272791 119869 272839 119897
rect 272529 119835 272839 119869
rect 272529 119807 272577 119835
rect 272605 119807 272639 119835
rect 272667 119807 272701 119835
rect 272729 119807 272763 119835
rect 272791 119807 272839 119835
rect 272529 119773 272839 119807
rect 272529 119745 272577 119773
rect 272605 119745 272639 119773
rect 272667 119745 272701 119773
rect 272729 119745 272763 119773
rect 272791 119745 272839 119773
rect 272529 110959 272839 119745
rect 272529 110931 272577 110959
rect 272605 110931 272639 110959
rect 272667 110931 272701 110959
rect 272729 110931 272763 110959
rect 272791 110931 272839 110959
rect 272529 110897 272839 110931
rect 272529 110869 272577 110897
rect 272605 110869 272639 110897
rect 272667 110869 272701 110897
rect 272729 110869 272763 110897
rect 272791 110869 272839 110897
rect 272529 110835 272839 110869
rect 272529 110807 272577 110835
rect 272605 110807 272639 110835
rect 272667 110807 272701 110835
rect 272729 110807 272763 110835
rect 272791 110807 272839 110835
rect 272529 110773 272839 110807
rect 272529 110745 272577 110773
rect 272605 110745 272639 110773
rect 272667 110745 272701 110773
rect 272729 110745 272763 110773
rect 272791 110745 272839 110773
rect 272529 101959 272839 110745
rect 272529 101931 272577 101959
rect 272605 101931 272639 101959
rect 272667 101931 272701 101959
rect 272729 101931 272763 101959
rect 272791 101931 272839 101959
rect 272529 101897 272839 101931
rect 272529 101869 272577 101897
rect 272605 101869 272639 101897
rect 272667 101869 272701 101897
rect 272729 101869 272763 101897
rect 272791 101869 272839 101897
rect 272529 101835 272839 101869
rect 272529 101807 272577 101835
rect 272605 101807 272639 101835
rect 272667 101807 272701 101835
rect 272729 101807 272763 101835
rect 272791 101807 272839 101835
rect 272529 101773 272839 101807
rect 272529 101745 272577 101773
rect 272605 101745 272639 101773
rect 272667 101745 272701 101773
rect 272729 101745 272763 101773
rect 272791 101745 272839 101773
rect 272529 92959 272839 101745
rect 272529 92931 272577 92959
rect 272605 92931 272639 92959
rect 272667 92931 272701 92959
rect 272729 92931 272763 92959
rect 272791 92931 272839 92959
rect 272529 92897 272839 92931
rect 272529 92869 272577 92897
rect 272605 92869 272639 92897
rect 272667 92869 272701 92897
rect 272729 92869 272763 92897
rect 272791 92869 272839 92897
rect 272529 92835 272839 92869
rect 272529 92807 272577 92835
rect 272605 92807 272639 92835
rect 272667 92807 272701 92835
rect 272729 92807 272763 92835
rect 272791 92807 272839 92835
rect 272529 92773 272839 92807
rect 272529 92745 272577 92773
rect 272605 92745 272639 92773
rect 272667 92745 272701 92773
rect 272729 92745 272763 92773
rect 272791 92745 272839 92773
rect 272529 83959 272839 92745
rect 272529 83931 272577 83959
rect 272605 83931 272639 83959
rect 272667 83931 272701 83959
rect 272729 83931 272763 83959
rect 272791 83931 272839 83959
rect 272529 83897 272839 83931
rect 272529 83869 272577 83897
rect 272605 83869 272639 83897
rect 272667 83869 272701 83897
rect 272729 83869 272763 83897
rect 272791 83869 272839 83897
rect 272529 83835 272839 83869
rect 272529 83807 272577 83835
rect 272605 83807 272639 83835
rect 272667 83807 272701 83835
rect 272729 83807 272763 83835
rect 272791 83807 272839 83835
rect 272529 83773 272839 83807
rect 272529 83745 272577 83773
rect 272605 83745 272639 83773
rect 272667 83745 272701 83773
rect 272729 83745 272763 83773
rect 272791 83745 272839 83773
rect 272529 74959 272839 83745
rect 272529 74931 272577 74959
rect 272605 74931 272639 74959
rect 272667 74931 272701 74959
rect 272729 74931 272763 74959
rect 272791 74931 272839 74959
rect 272529 74897 272839 74931
rect 272529 74869 272577 74897
rect 272605 74869 272639 74897
rect 272667 74869 272701 74897
rect 272729 74869 272763 74897
rect 272791 74869 272839 74897
rect 272529 74835 272839 74869
rect 272529 74807 272577 74835
rect 272605 74807 272639 74835
rect 272667 74807 272701 74835
rect 272729 74807 272763 74835
rect 272791 74807 272839 74835
rect 272529 74773 272839 74807
rect 272529 74745 272577 74773
rect 272605 74745 272639 74773
rect 272667 74745 272701 74773
rect 272729 74745 272763 74773
rect 272791 74745 272839 74773
rect 272529 65959 272839 74745
rect 272529 65931 272577 65959
rect 272605 65931 272639 65959
rect 272667 65931 272701 65959
rect 272729 65931 272763 65959
rect 272791 65931 272839 65959
rect 272529 65897 272839 65931
rect 272529 65869 272577 65897
rect 272605 65869 272639 65897
rect 272667 65869 272701 65897
rect 272729 65869 272763 65897
rect 272791 65869 272839 65897
rect 272529 65835 272839 65869
rect 272529 65807 272577 65835
rect 272605 65807 272639 65835
rect 272667 65807 272701 65835
rect 272729 65807 272763 65835
rect 272791 65807 272839 65835
rect 272529 65773 272839 65807
rect 272529 65745 272577 65773
rect 272605 65745 272639 65773
rect 272667 65745 272701 65773
rect 272729 65745 272763 65773
rect 272791 65745 272839 65773
rect 272529 56959 272839 65745
rect 272529 56931 272577 56959
rect 272605 56931 272639 56959
rect 272667 56931 272701 56959
rect 272729 56931 272763 56959
rect 272791 56931 272839 56959
rect 272529 56897 272839 56931
rect 272529 56869 272577 56897
rect 272605 56869 272639 56897
rect 272667 56869 272701 56897
rect 272729 56869 272763 56897
rect 272791 56869 272839 56897
rect 272529 56835 272839 56869
rect 272529 56807 272577 56835
rect 272605 56807 272639 56835
rect 272667 56807 272701 56835
rect 272729 56807 272763 56835
rect 272791 56807 272839 56835
rect 272529 56773 272839 56807
rect 272529 56745 272577 56773
rect 272605 56745 272639 56773
rect 272667 56745 272701 56773
rect 272729 56745 272763 56773
rect 272791 56745 272839 56773
rect 272529 47959 272839 56745
rect 272529 47931 272577 47959
rect 272605 47931 272639 47959
rect 272667 47931 272701 47959
rect 272729 47931 272763 47959
rect 272791 47931 272839 47959
rect 272529 47897 272839 47931
rect 272529 47869 272577 47897
rect 272605 47869 272639 47897
rect 272667 47869 272701 47897
rect 272729 47869 272763 47897
rect 272791 47869 272839 47897
rect 272529 47835 272839 47869
rect 272529 47807 272577 47835
rect 272605 47807 272639 47835
rect 272667 47807 272701 47835
rect 272729 47807 272763 47835
rect 272791 47807 272839 47835
rect 272529 47773 272839 47807
rect 272529 47745 272577 47773
rect 272605 47745 272639 47773
rect 272667 47745 272701 47773
rect 272729 47745 272763 47773
rect 272791 47745 272839 47773
rect 272529 38959 272839 47745
rect 272529 38931 272577 38959
rect 272605 38931 272639 38959
rect 272667 38931 272701 38959
rect 272729 38931 272763 38959
rect 272791 38931 272839 38959
rect 272529 38897 272839 38931
rect 272529 38869 272577 38897
rect 272605 38869 272639 38897
rect 272667 38869 272701 38897
rect 272729 38869 272763 38897
rect 272791 38869 272839 38897
rect 272529 38835 272839 38869
rect 272529 38807 272577 38835
rect 272605 38807 272639 38835
rect 272667 38807 272701 38835
rect 272729 38807 272763 38835
rect 272791 38807 272839 38835
rect 272529 38773 272839 38807
rect 272529 38745 272577 38773
rect 272605 38745 272639 38773
rect 272667 38745 272701 38773
rect 272729 38745 272763 38773
rect 272791 38745 272839 38773
rect 272529 29959 272839 38745
rect 272529 29931 272577 29959
rect 272605 29931 272639 29959
rect 272667 29931 272701 29959
rect 272729 29931 272763 29959
rect 272791 29931 272839 29959
rect 272529 29897 272839 29931
rect 272529 29869 272577 29897
rect 272605 29869 272639 29897
rect 272667 29869 272701 29897
rect 272729 29869 272763 29897
rect 272791 29869 272839 29897
rect 272529 29835 272839 29869
rect 272529 29807 272577 29835
rect 272605 29807 272639 29835
rect 272667 29807 272701 29835
rect 272729 29807 272763 29835
rect 272791 29807 272839 29835
rect 272529 29773 272839 29807
rect 272529 29745 272577 29773
rect 272605 29745 272639 29773
rect 272667 29745 272701 29773
rect 272729 29745 272763 29773
rect 272791 29745 272839 29773
rect 272529 20959 272839 29745
rect 272529 20931 272577 20959
rect 272605 20931 272639 20959
rect 272667 20931 272701 20959
rect 272729 20931 272763 20959
rect 272791 20931 272839 20959
rect 272529 20897 272839 20931
rect 272529 20869 272577 20897
rect 272605 20869 272639 20897
rect 272667 20869 272701 20897
rect 272729 20869 272763 20897
rect 272791 20869 272839 20897
rect 272529 20835 272839 20869
rect 272529 20807 272577 20835
rect 272605 20807 272639 20835
rect 272667 20807 272701 20835
rect 272729 20807 272763 20835
rect 272791 20807 272839 20835
rect 272529 20773 272839 20807
rect 272529 20745 272577 20773
rect 272605 20745 272639 20773
rect 272667 20745 272701 20773
rect 272729 20745 272763 20773
rect 272791 20745 272839 20773
rect 272529 11959 272839 20745
rect 272529 11931 272577 11959
rect 272605 11931 272639 11959
rect 272667 11931 272701 11959
rect 272729 11931 272763 11959
rect 272791 11931 272839 11959
rect 272529 11897 272839 11931
rect 272529 11869 272577 11897
rect 272605 11869 272639 11897
rect 272667 11869 272701 11897
rect 272729 11869 272763 11897
rect 272791 11869 272839 11897
rect 272529 11835 272839 11869
rect 272529 11807 272577 11835
rect 272605 11807 272639 11835
rect 272667 11807 272701 11835
rect 272729 11807 272763 11835
rect 272791 11807 272839 11835
rect 272529 11773 272839 11807
rect 272529 11745 272577 11773
rect 272605 11745 272639 11773
rect 272667 11745 272701 11773
rect 272729 11745 272763 11773
rect 272791 11745 272839 11773
rect 272529 2959 272839 11745
rect 272529 2931 272577 2959
rect 272605 2931 272639 2959
rect 272667 2931 272701 2959
rect 272729 2931 272763 2959
rect 272791 2931 272839 2959
rect 272529 2897 272839 2931
rect 272529 2869 272577 2897
rect 272605 2869 272639 2897
rect 272667 2869 272701 2897
rect 272729 2869 272763 2897
rect 272791 2869 272839 2897
rect 272529 2835 272839 2869
rect 272529 2807 272577 2835
rect 272605 2807 272639 2835
rect 272667 2807 272701 2835
rect 272729 2807 272763 2835
rect 272791 2807 272839 2835
rect 272529 2773 272839 2807
rect 272529 2745 272577 2773
rect 272605 2745 272639 2773
rect 272667 2745 272701 2773
rect 272729 2745 272763 2773
rect 272791 2745 272839 2773
rect 272529 904 272839 2745
rect 272529 876 272577 904
rect 272605 876 272639 904
rect 272667 876 272701 904
rect 272729 876 272763 904
rect 272791 876 272839 904
rect 272529 842 272839 876
rect 272529 814 272577 842
rect 272605 814 272639 842
rect 272667 814 272701 842
rect 272729 814 272763 842
rect 272791 814 272839 842
rect 272529 780 272839 814
rect 272529 752 272577 780
rect 272605 752 272639 780
rect 272667 752 272701 780
rect 272729 752 272763 780
rect 272791 752 272839 780
rect 272529 718 272839 752
rect 272529 690 272577 718
rect 272605 690 272639 718
rect 272667 690 272701 718
rect 272729 690 272763 718
rect 272791 690 272839 718
rect 272529 162 272839 690
rect 274389 299670 274699 299718
rect 274389 299642 274437 299670
rect 274465 299642 274499 299670
rect 274527 299642 274561 299670
rect 274589 299642 274623 299670
rect 274651 299642 274699 299670
rect 274389 299608 274699 299642
rect 274389 299580 274437 299608
rect 274465 299580 274499 299608
rect 274527 299580 274561 299608
rect 274589 299580 274623 299608
rect 274651 299580 274699 299608
rect 274389 299546 274699 299580
rect 274389 299518 274437 299546
rect 274465 299518 274499 299546
rect 274527 299518 274561 299546
rect 274589 299518 274623 299546
rect 274651 299518 274699 299546
rect 274389 299484 274699 299518
rect 274389 299456 274437 299484
rect 274465 299456 274499 299484
rect 274527 299456 274561 299484
rect 274589 299456 274623 299484
rect 274651 299456 274699 299484
rect 274389 293959 274699 299456
rect 274389 293931 274437 293959
rect 274465 293931 274499 293959
rect 274527 293931 274561 293959
rect 274589 293931 274623 293959
rect 274651 293931 274699 293959
rect 274389 293897 274699 293931
rect 274389 293869 274437 293897
rect 274465 293869 274499 293897
rect 274527 293869 274561 293897
rect 274589 293869 274623 293897
rect 274651 293869 274699 293897
rect 274389 293835 274699 293869
rect 274389 293807 274437 293835
rect 274465 293807 274499 293835
rect 274527 293807 274561 293835
rect 274589 293807 274623 293835
rect 274651 293807 274699 293835
rect 274389 293773 274699 293807
rect 274389 293745 274437 293773
rect 274465 293745 274499 293773
rect 274527 293745 274561 293773
rect 274589 293745 274623 293773
rect 274651 293745 274699 293773
rect 274389 284959 274699 293745
rect 274389 284931 274437 284959
rect 274465 284931 274499 284959
rect 274527 284931 274561 284959
rect 274589 284931 274623 284959
rect 274651 284931 274699 284959
rect 274389 284897 274699 284931
rect 274389 284869 274437 284897
rect 274465 284869 274499 284897
rect 274527 284869 274561 284897
rect 274589 284869 274623 284897
rect 274651 284869 274699 284897
rect 274389 284835 274699 284869
rect 274389 284807 274437 284835
rect 274465 284807 274499 284835
rect 274527 284807 274561 284835
rect 274589 284807 274623 284835
rect 274651 284807 274699 284835
rect 274389 284773 274699 284807
rect 274389 284745 274437 284773
rect 274465 284745 274499 284773
rect 274527 284745 274561 284773
rect 274589 284745 274623 284773
rect 274651 284745 274699 284773
rect 274389 275959 274699 284745
rect 274389 275931 274437 275959
rect 274465 275931 274499 275959
rect 274527 275931 274561 275959
rect 274589 275931 274623 275959
rect 274651 275931 274699 275959
rect 274389 275897 274699 275931
rect 274389 275869 274437 275897
rect 274465 275869 274499 275897
rect 274527 275869 274561 275897
rect 274589 275869 274623 275897
rect 274651 275869 274699 275897
rect 274389 275835 274699 275869
rect 274389 275807 274437 275835
rect 274465 275807 274499 275835
rect 274527 275807 274561 275835
rect 274589 275807 274623 275835
rect 274651 275807 274699 275835
rect 274389 275773 274699 275807
rect 274389 275745 274437 275773
rect 274465 275745 274499 275773
rect 274527 275745 274561 275773
rect 274589 275745 274623 275773
rect 274651 275745 274699 275773
rect 274389 266959 274699 275745
rect 274389 266931 274437 266959
rect 274465 266931 274499 266959
rect 274527 266931 274561 266959
rect 274589 266931 274623 266959
rect 274651 266931 274699 266959
rect 274389 266897 274699 266931
rect 274389 266869 274437 266897
rect 274465 266869 274499 266897
rect 274527 266869 274561 266897
rect 274589 266869 274623 266897
rect 274651 266869 274699 266897
rect 274389 266835 274699 266869
rect 274389 266807 274437 266835
rect 274465 266807 274499 266835
rect 274527 266807 274561 266835
rect 274589 266807 274623 266835
rect 274651 266807 274699 266835
rect 274389 266773 274699 266807
rect 274389 266745 274437 266773
rect 274465 266745 274499 266773
rect 274527 266745 274561 266773
rect 274589 266745 274623 266773
rect 274651 266745 274699 266773
rect 274389 257959 274699 266745
rect 274389 257931 274437 257959
rect 274465 257931 274499 257959
rect 274527 257931 274561 257959
rect 274589 257931 274623 257959
rect 274651 257931 274699 257959
rect 274389 257897 274699 257931
rect 274389 257869 274437 257897
rect 274465 257869 274499 257897
rect 274527 257869 274561 257897
rect 274589 257869 274623 257897
rect 274651 257869 274699 257897
rect 274389 257835 274699 257869
rect 274389 257807 274437 257835
rect 274465 257807 274499 257835
rect 274527 257807 274561 257835
rect 274589 257807 274623 257835
rect 274651 257807 274699 257835
rect 274389 257773 274699 257807
rect 274389 257745 274437 257773
rect 274465 257745 274499 257773
rect 274527 257745 274561 257773
rect 274589 257745 274623 257773
rect 274651 257745 274699 257773
rect 274389 248959 274699 257745
rect 274389 248931 274437 248959
rect 274465 248931 274499 248959
rect 274527 248931 274561 248959
rect 274589 248931 274623 248959
rect 274651 248931 274699 248959
rect 274389 248897 274699 248931
rect 274389 248869 274437 248897
rect 274465 248869 274499 248897
rect 274527 248869 274561 248897
rect 274589 248869 274623 248897
rect 274651 248869 274699 248897
rect 274389 248835 274699 248869
rect 274389 248807 274437 248835
rect 274465 248807 274499 248835
rect 274527 248807 274561 248835
rect 274589 248807 274623 248835
rect 274651 248807 274699 248835
rect 274389 248773 274699 248807
rect 274389 248745 274437 248773
rect 274465 248745 274499 248773
rect 274527 248745 274561 248773
rect 274589 248745 274623 248773
rect 274651 248745 274699 248773
rect 274389 239959 274699 248745
rect 274389 239931 274437 239959
rect 274465 239931 274499 239959
rect 274527 239931 274561 239959
rect 274589 239931 274623 239959
rect 274651 239931 274699 239959
rect 274389 239897 274699 239931
rect 274389 239869 274437 239897
rect 274465 239869 274499 239897
rect 274527 239869 274561 239897
rect 274589 239869 274623 239897
rect 274651 239869 274699 239897
rect 274389 239835 274699 239869
rect 274389 239807 274437 239835
rect 274465 239807 274499 239835
rect 274527 239807 274561 239835
rect 274589 239807 274623 239835
rect 274651 239807 274699 239835
rect 274389 239773 274699 239807
rect 274389 239745 274437 239773
rect 274465 239745 274499 239773
rect 274527 239745 274561 239773
rect 274589 239745 274623 239773
rect 274651 239745 274699 239773
rect 274389 230959 274699 239745
rect 274389 230931 274437 230959
rect 274465 230931 274499 230959
rect 274527 230931 274561 230959
rect 274589 230931 274623 230959
rect 274651 230931 274699 230959
rect 274389 230897 274699 230931
rect 274389 230869 274437 230897
rect 274465 230869 274499 230897
rect 274527 230869 274561 230897
rect 274589 230869 274623 230897
rect 274651 230869 274699 230897
rect 274389 230835 274699 230869
rect 274389 230807 274437 230835
rect 274465 230807 274499 230835
rect 274527 230807 274561 230835
rect 274589 230807 274623 230835
rect 274651 230807 274699 230835
rect 274389 230773 274699 230807
rect 274389 230745 274437 230773
rect 274465 230745 274499 230773
rect 274527 230745 274561 230773
rect 274589 230745 274623 230773
rect 274651 230745 274699 230773
rect 274389 221959 274699 230745
rect 274389 221931 274437 221959
rect 274465 221931 274499 221959
rect 274527 221931 274561 221959
rect 274589 221931 274623 221959
rect 274651 221931 274699 221959
rect 274389 221897 274699 221931
rect 274389 221869 274437 221897
rect 274465 221869 274499 221897
rect 274527 221869 274561 221897
rect 274589 221869 274623 221897
rect 274651 221869 274699 221897
rect 274389 221835 274699 221869
rect 274389 221807 274437 221835
rect 274465 221807 274499 221835
rect 274527 221807 274561 221835
rect 274589 221807 274623 221835
rect 274651 221807 274699 221835
rect 274389 221773 274699 221807
rect 274389 221745 274437 221773
rect 274465 221745 274499 221773
rect 274527 221745 274561 221773
rect 274589 221745 274623 221773
rect 274651 221745 274699 221773
rect 274389 212959 274699 221745
rect 274389 212931 274437 212959
rect 274465 212931 274499 212959
rect 274527 212931 274561 212959
rect 274589 212931 274623 212959
rect 274651 212931 274699 212959
rect 274389 212897 274699 212931
rect 274389 212869 274437 212897
rect 274465 212869 274499 212897
rect 274527 212869 274561 212897
rect 274589 212869 274623 212897
rect 274651 212869 274699 212897
rect 274389 212835 274699 212869
rect 274389 212807 274437 212835
rect 274465 212807 274499 212835
rect 274527 212807 274561 212835
rect 274589 212807 274623 212835
rect 274651 212807 274699 212835
rect 274389 212773 274699 212807
rect 274389 212745 274437 212773
rect 274465 212745 274499 212773
rect 274527 212745 274561 212773
rect 274589 212745 274623 212773
rect 274651 212745 274699 212773
rect 274389 203959 274699 212745
rect 274389 203931 274437 203959
rect 274465 203931 274499 203959
rect 274527 203931 274561 203959
rect 274589 203931 274623 203959
rect 274651 203931 274699 203959
rect 274389 203897 274699 203931
rect 274389 203869 274437 203897
rect 274465 203869 274499 203897
rect 274527 203869 274561 203897
rect 274589 203869 274623 203897
rect 274651 203869 274699 203897
rect 274389 203835 274699 203869
rect 274389 203807 274437 203835
rect 274465 203807 274499 203835
rect 274527 203807 274561 203835
rect 274589 203807 274623 203835
rect 274651 203807 274699 203835
rect 274389 203773 274699 203807
rect 274389 203745 274437 203773
rect 274465 203745 274499 203773
rect 274527 203745 274561 203773
rect 274589 203745 274623 203773
rect 274651 203745 274699 203773
rect 274389 194959 274699 203745
rect 274389 194931 274437 194959
rect 274465 194931 274499 194959
rect 274527 194931 274561 194959
rect 274589 194931 274623 194959
rect 274651 194931 274699 194959
rect 274389 194897 274699 194931
rect 274389 194869 274437 194897
rect 274465 194869 274499 194897
rect 274527 194869 274561 194897
rect 274589 194869 274623 194897
rect 274651 194869 274699 194897
rect 274389 194835 274699 194869
rect 274389 194807 274437 194835
rect 274465 194807 274499 194835
rect 274527 194807 274561 194835
rect 274589 194807 274623 194835
rect 274651 194807 274699 194835
rect 274389 194773 274699 194807
rect 274389 194745 274437 194773
rect 274465 194745 274499 194773
rect 274527 194745 274561 194773
rect 274589 194745 274623 194773
rect 274651 194745 274699 194773
rect 274389 185959 274699 194745
rect 274389 185931 274437 185959
rect 274465 185931 274499 185959
rect 274527 185931 274561 185959
rect 274589 185931 274623 185959
rect 274651 185931 274699 185959
rect 274389 185897 274699 185931
rect 274389 185869 274437 185897
rect 274465 185869 274499 185897
rect 274527 185869 274561 185897
rect 274589 185869 274623 185897
rect 274651 185869 274699 185897
rect 274389 185835 274699 185869
rect 274389 185807 274437 185835
rect 274465 185807 274499 185835
rect 274527 185807 274561 185835
rect 274589 185807 274623 185835
rect 274651 185807 274699 185835
rect 274389 185773 274699 185807
rect 274389 185745 274437 185773
rect 274465 185745 274499 185773
rect 274527 185745 274561 185773
rect 274589 185745 274623 185773
rect 274651 185745 274699 185773
rect 274389 176959 274699 185745
rect 274389 176931 274437 176959
rect 274465 176931 274499 176959
rect 274527 176931 274561 176959
rect 274589 176931 274623 176959
rect 274651 176931 274699 176959
rect 274389 176897 274699 176931
rect 274389 176869 274437 176897
rect 274465 176869 274499 176897
rect 274527 176869 274561 176897
rect 274589 176869 274623 176897
rect 274651 176869 274699 176897
rect 274389 176835 274699 176869
rect 274389 176807 274437 176835
rect 274465 176807 274499 176835
rect 274527 176807 274561 176835
rect 274589 176807 274623 176835
rect 274651 176807 274699 176835
rect 274389 176773 274699 176807
rect 274389 176745 274437 176773
rect 274465 176745 274499 176773
rect 274527 176745 274561 176773
rect 274589 176745 274623 176773
rect 274651 176745 274699 176773
rect 274389 167959 274699 176745
rect 274389 167931 274437 167959
rect 274465 167931 274499 167959
rect 274527 167931 274561 167959
rect 274589 167931 274623 167959
rect 274651 167931 274699 167959
rect 274389 167897 274699 167931
rect 274389 167869 274437 167897
rect 274465 167869 274499 167897
rect 274527 167869 274561 167897
rect 274589 167869 274623 167897
rect 274651 167869 274699 167897
rect 274389 167835 274699 167869
rect 274389 167807 274437 167835
rect 274465 167807 274499 167835
rect 274527 167807 274561 167835
rect 274589 167807 274623 167835
rect 274651 167807 274699 167835
rect 274389 167773 274699 167807
rect 274389 167745 274437 167773
rect 274465 167745 274499 167773
rect 274527 167745 274561 167773
rect 274589 167745 274623 167773
rect 274651 167745 274699 167773
rect 274389 158959 274699 167745
rect 274389 158931 274437 158959
rect 274465 158931 274499 158959
rect 274527 158931 274561 158959
rect 274589 158931 274623 158959
rect 274651 158931 274699 158959
rect 274389 158897 274699 158931
rect 274389 158869 274437 158897
rect 274465 158869 274499 158897
rect 274527 158869 274561 158897
rect 274589 158869 274623 158897
rect 274651 158869 274699 158897
rect 274389 158835 274699 158869
rect 274389 158807 274437 158835
rect 274465 158807 274499 158835
rect 274527 158807 274561 158835
rect 274589 158807 274623 158835
rect 274651 158807 274699 158835
rect 274389 158773 274699 158807
rect 274389 158745 274437 158773
rect 274465 158745 274499 158773
rect 274527 158745 274561 158773
rect 274589 158745 274623 158773
rect 274651 158745 274699 158773
rect 274389 149959 274699 158745
rect 274389 149931 274437 149959
rect 274465 149931 274499 149959
rect 274527 149931 274561 149959
rect 274589 149931 274623 149959
rect 274651 149931 274699 149959
rect 274389 149897 274699 149931
rect 274389 149869 274437 149897
rect 274465 149869 274499 149897
rect 274527 149869 274561 149897
rect 274589 149869 274623 149897
rect 274651 149869 274699 149897
rect 274389 149835 274699 149869
rect 274389 149807 274437 149835
rect 274465 149807 274499 149835
rect 274527 149807 274561 149835
rect 274589 149807 274623 149835
rect 274651 149807 274699 149835
rect 274389 149773 274699 149807
rect 274389 149745 274437 149773
rect 274465 149745 274499 149773
rect 274527 149745 274561 149773
rect 274589 149745 274623 149773
rect 274651 149745 274699 149773
rect 274389 140959 274699 149745
rect 274389 140931 274437 140959
rect 274465 140931 274499 140959
rect 274527 140931 274561 140959
rect 274589 140931 274623 140959
rect 274651 140931 274699 140959
rect 274389 140897 274699 140931
rect 274389 140869 274437 140897
rect 274465 140869 274499 140897
rect 274527 140869 274561 140897
rect 274589 140869 274623 140897
rect 274651 140869 274699 140897
rect 274389 140835 274699 140869
rect 274389 140807 274437 140835
rect 274465 140807 274499 140835
rect 274527 140807 274561 140835
rect 274589 140807 274623 140835
rect 274651 140807 274699 140835
rect 274389 140773 274699 140807
rect 274389 140745 274437 140773
rect 274465 140745 274499 140773
rect 274527 140745 274561 140773
rect 274589 140745 274623 140773
rect 274651 140745 274699 140773
rect 274389 131959 274699 140745
rect 274389 131931 274437 131959
rect 274465 131931 274499 131959
rect 274527 131931 274561 131959
rect 274589 131931 274623 131959
rect 274651 131931 274699 131959
rect 274389 131897 274699 131931
rect 274389 131869 274437 131897
rect 274465 131869 274499 131897
rect 274527 131869 274561 131897
rect 274589 131869 274623 131897
rect 274651 131869 274699 131897
rect 274389 131835 274699 131869
rect 274389 131807 274437 131835
rect 274465 131807 274499 131835
rect 274527 131807 274561 131835
rect 274589 131807 274623 131835
rect 274651 131807 274699 131835
rect 274389 131773 274699 131807
rect 274389 131745 274437 131773
rect 274465 131745 274499 131773
rect 274527 131745 274561 131773
rect 274589 131745 274623 131773
rect 274651 131745 274699 131773
rect 274389 122959 274699 131745
rect 274389 122931 274437 122959
rect 274465 122931 274499 122959
rect 274527 122931 274561 122959
rect 274589 122931 274623 122959
rect 274651 122931 274699 122959
rect 274389 122897 274699 122931
rect 274389 122869 274437 122897
rect 274465 122869 274499 122897
rect 274527 122869 274561 122897
rect 274589 122869 274623 122897
rect 274651 122869 274699 122897
rect 274389 122835 274699 122869
rect 274389 122807 274437 122835
rect 274465 122807 274499 122835
rect 274527 122807 274561 122835
rect 274589 122807 274623 122835
rect 274651 122807 274699 122835
rect 274389 122773 274699 122807
rect 274389 122745 274437 122773
rect 274465 122745 274499 122773
rect 274527 122745 274561 122773
rect 274589 122745 274623 122773
rect 274651 122745 274699 122773
rect 274389 113959 274699 122745
rect 274389 113931 274437 113959
rect 274465 113931 274499 113959
rect 274527 113931 274561 113959
rect 274589 113931 274623 113959
rect 274651 113931 274699 113959
rect 274389 113897 274699 113931
rect 274389 113869 274437 113897
rect 274465 113869 274499 113897
rect 274527 113869 274561 113897
rect 274589 113869 274623 113897
rect 274651 113869 274699 113897
rect 274389 113835 274699 113869
rect 274389 113807 274437 113835
rect 274465 113807 274499 113835
rect 274527 113807 274561 113835
rect 274589 113807 274623 113835
rect 274651 113807 274699 113835
rect 274389 113773 274699 113807
rect 274389 113745 274437 113773
rect 274465 113745 274499 113773
rect 274527 113745 274561 113773
rect 274589 113745 274623 113773
rect 274651 113745 274699 113773
rect 274389 104959 274699 113745
rect 274389 104931 274437 104959
rect 274465 104931 274499 104959
rect 274527 104931 274561 104959
rect 274589 104931 274623 104959
rect 274651 104931 274699 104959
rect 274389 104897 274699 104931
rect 274389 104869 274437 104897
rect 274465 104869 274499 104897
rect 274527 104869 274561 104897
rect 274589 104869 274623 104897
rect 274651 104869 274699 104897
rect 274389 104835 274699 104869
rect 274389 104807 274437 104835
rect 274465 104807 274499 104835
rect 274527 104807 274561 104835
rect 274589 104807 274623 104835
rect 274651 104807 274699 104835
rect 274389 104773 274699 104807
rect 274389 104745 274437 104773
rect 274465 104745 274499 104773
rect 274527 104745 274561 104773
rect 274589 104745 274623 104773
rect 274651 104745 274699 104773
rect 274389 95959 274699 104745
rect 274389 95931 274437 95959
rect 274465 95931 274499 95959
rect 274527 95931 274561 95959
rect 274589 95931 274623 95959
rect 274651 95931 274699 95959
rect 274389 95897 274699 95931
rect 274389 95869 274437 95897
rect 274465 95869 274499 95897
rect 274527 95869 274561 95897
rect 274589 95869 274623 95897
rect 274651 95869 274699 95897
rect 274389 95835 274699 95869
rect 274389 95807 274437 95835
rect 274465 95807 274499 95835
rect 274527 95807 274561 95835
rect 274589 95807 274623 95835
rect 274651 95807 274699 95835
rect 274389 95773 274699 95807
rect 274389 95745 274437 95773
rect 274465 95745 274499 95773
rect 274527 95745 274561 95773
rect 274589 95745 274623 95773
rect 274651 95745 274699 95773
rect 274389 86959 274699 95745
rect 274389 86931 274437 86959
rect 274465 86931 274499 86959
rect 274527 86931 274561 86959
rect 274589 86931 274623 86959
rect 274651 86931 274699 86959
rect 274389 86897 274699 86931
rect 274389 86869 274437 86897
rect 274465 86869 274499 86897
rect 274527 86869 274561 86897
rect 274589 86869 274623 86897
rect 274651 86869 274699 86897
rect 274389 86835 274699 86869
rect 274389 86807 274437 86835
rect 274465 86807 274499 86835
rect 274527 86807 274561 86835
rect 274589 86807 274623 86835
rect 274651 86807 274699 86835
rect 274389 86773 274699 86807
rect 274389 86745 274437 86773
rect 274465 86745 274499 86773
rect 274527 86745 274561 86773
rect 274589 86745 274623 86773
rect 274651 86745 274699 86773
rect 274389 77959 274699 86745
rect 274389 77931 274437 77959
rect 274465 77931 274499 77959
rect 274527 77931 274561 77959
rect 274589 77931 274623 77959
rect 274651 77931 274699 77959
rect 274389 77897 274699 77931
rect 274389 77869 274437 77897
rect 274465 77869 274499 77897
rect 274527 77869 274561 77897
rect 274589 77869 274623 77897
rect 274651 77869 274699 77897
rect 274389 77835 274699 77869
rect 274389 77807 274437 77835
rect 274465 77807 274499 77835
rect 274527 77807 274561 77835
rect 274589 77807 274623 77835
rect 274651 77807 274699 77835
rect 274389 77773 274699 77807
rect 274389 77745 274437 77773
rect 274465 77745 274499 77773
rect 274527 77745 274561 77773
rect 274589 77745 274623 77773
rect 274651 77745 274699 77773
rect 274389 68959 274699 77745
rect 274389 68931 274437 68959
rect 274465 68931 274499 68959
rect 274527 68931 274561 68959
rect 274589 68931 274623 68959
rect 274651 68931 274699 68959
rect 274389 68897 274699 68931
rect 274389 68869 274437 68897
rect 274465 68869 274499 68897
rect 274527 68869 274561 68897
rect 274589 68869 274623 68897
rect 274651 68869 274699 68897
rect 274389 68835 274699 68869
rect 274389 68807 274437 68835
rect 274465 68807 274499 68835
rect 274527 68807 274561 68835
rect 274589 68807 274623 68835
rect 274651 68807 274699 68835
rect 274389 68773 274699 68807
rect 274389 68745 274437 68773
rect 274465 68745 274499 68773
rect 274527 68745 274561 68773
rect 274589 68745 274623 68773
rect 274651 68745 274699 68773
rect 274389 59959 274699 68745
rect 274389 59931 274437 59959
rect 274465 59931 274499 59959
rect 274527 59931 274561 59959
rect 274589 59931 274623 59959
rect 274651 59931 274699 59959
rect 274389 59897 274699 59931
rect 274389 59869 274437 59897
rect 274465 59869 274499 59897
rect 274527 59869 274561 59897
rect 274589 59869 274623 59897
rect 274651 59869 274699 59897
rect 274389 59835 274699 59869
rect 274389 59807 274437 59835
rect 274465 59807 274499 59835
rect 274527 59807 274561 59835
rect 274589 59807 274623 59835
rect 274651 59807 274699 59835
rect 274389 59773 274699 59807
rect 274389 59745 274437 59773
rect 274465 59745 274499 59773
rect 274527 59745 274561 59773
rect 274589 59745 274623 59773
rect 274651 59745 274699 59773
rect 274389 50959 274699 59745
rect 274389 50931 274437 50959
rect 274465 50931 274499 50959
rect 274527 50931 274561 50959
rect 274589 50931 274623 50959
rect 274651 50931 274699 50959
rect 274389 50897 274699 50931
rect 274389 50869 274437 50897
rect 274465 50869 274499 50897
rect 274527 50869 274561 50897
rect 274589 50869 274623 50897
rect 274651 50869 274699 50897
rect 274389 50835 274699 50869
rect 274389 50807 274437 50835
rect 274465 50807 274499 50835
rect 274527 50807 274561 50835
rect 274589 50807 274623 50835
rect 274651 50807 274699 50835
rect 274389 50773 274699 50807
rect 274389 50745 274437 50773
rect 274465 50745 274499 50773
rect 274527 50745 274561 50773
rect 274589 50745 274623 50773
rect 274651 50745 274699 50773
rect 274389 41959 274699 50745
rect 274389 41931 274437 41959
rect 274465 41931 274499 41959
rect 274527 41931 274561 41959
rect 274589 41931 274623 41959
rect 274651 41931 274699 41959
rect 274389 41897 274699 41931
rect 274389 41869 274437 41897
rect 274465 41869 274499 41897
rect 274527 41869 274561 41897
rect 274589 41869 274623 41897
rect 274651 41869 274699 41897
rect 274389 41835 274699 41869
rect 274389 41807 274437 41835
rect 274465 41807 274499 41835
rect 274527 41807 274561 41835
rect 274589 41807 274623 41835
rect 274651 41807 274699 41835
rect 274389 41773 274699 41807
rect 274389 41745 274437 41773
rect 274465 41745 274499 41773
rect 274527 41745 274561 41773
rect 274589 41745 274623 41773
rect 274651 41745 274699 41773
rect 274389 32959 274699 41745
rect 274389 32931 274437 32959
rect 274465 32931 274499 32959
rect 274527 32931 274561 32959
rect 274589 32931 274623 32959
rect 274651 32931 274699 32959
rect 274389 32897 274699 32931
rect 274389 32869 274437 32897
rect 274465 32869 274499 32897
rect 274527 32869 274561 32897
rect 274589 32869 274623 32897
rect 274651 32869 274699 32897
rect 274389 32835 274699 32869
rect 274389 32807 274437 32835
rect 274465 32807 274499 32835
rect 274527 32807 274561 32835
rect 274589 32807 274623 32835
rect 274651 32807 274699 32835
rect 274389 32773 274699 32807
rect 274389 32745 274437 32773
rect 274465 32745 274499 32773
rect 274527 32745 274561 32773
rect 274589 32745 274623 32773
rect 274651 32745 274699 32773
rect 274389 23959 274699 32745
rect 274389 23931 274437 23959
rect 274465 23931 274499 23959
rect 274527 23931 274561 23959
rect 274589 23931 274623 23959
rect 274651 23931 274699 23959
rect 274389 23897 274699 23931
rect 274389 23869 274437 23897
rect 274465 23869 274499 23897
rect 274527 23869 274561 23897
rect 274589 23869 274623 23897
rect 274651 23869 274699 23897
rect 274389 23835 274699 23869
rect 274389 23807 274437 23835
rect 274465 23807 274499 23835
rect 274527 23807 274561 23835
rect 274589 23807 274623 23835
rect 274651 23807 274699 23835
rect 274389 23773 274699 23807
rect 274389 23745 274437 23773
rect 274465 23745 274499 23773
rect 274527 23745 274561 23773
rect 274589 23745 274623 23773
rect 274651 23745 274699 23773
rect 274389 14959 274699 23745
rect 274389 14931 274437 14959
rect 274465 14931 274499 14959
rect 274527 14931 274561 14959
rect 274589 14931 274623 14959
rect 274651 14931 274699 14959
rect 274389 14897 274699 14931
rect 274389 14869 274437 14897
rect 274465 14869 274499 14897
rect 274527 14869 274561 14897
rect 274589 14869 274623 14897
rect 274651 14869 274699 14897
rect 274389 14835 274699 14869
rect 274389 14807 274437 14835
rect 274465 14807 274499 14835
rect 274527 14807 274561 14835
rect 274589 14807 274623 14835
rect 274651 14807 274699 14835
rect 274389 14773 274699 14807
rect 274389 14745 274437 14773
rect 274465 14745 274499 14773
rect 274527 14745 274561 14773
rect 274589 14745 274623 14773
rect 274651 14745 274699 14773
rect 274389 5959 274699 14745
rect 274389 5931 274437 5959
rect 274465 5931 274499 5959
rect 274527 5931 274561 5959
rect 274589 5931 274623 5959
rect 274651 5931 274699 5959
rect 274389 5897 274699 5931
rect 274389 5869 274437 5897
rect 274465 5869 274499 5897
rect 274527 5869 274561 5897
rect 274589 5869 274623 5897
rect 274651 5869 274699 5897
rect 274389 5835 274699 5869
rect 274389 5807 274437 5835
rect 274465 5807 274499 5835
rect 274527 5807 274561 5835
rect 274589 5807 274623 5835
rect 274651 5807 274699 5835
rect 274389 5773 274699 5807
rect 274389 5745 274437 5773
rect 274465 5745 274499 5773
rect 274527 5745 274561 5773
rect 274589 5745 274623 5773
rect 274651 5745 274699 5773
rect 274389 424 274699 5745
rect 274389 396 274437 424
rect 274465 396 274499 424
rect 274527 396 274561 424
rect 274589 396 274623 424
rect 274651 396 274699 424
rect 274389 362 274699 396
rect 274389 334 274437 362
rect 274465 334 274499 362
rect 274527 334 274561 362
rect 274589 334 274623 362
rect 274651 334 274699 362
rect 274389 300 274699 334
rect 274389 272 274437 300
rect 274465 272 274499 300
rect 274527 272 274561 300
rect 274589 272 274623 300
rect 274651 272 274699 300
rect 274389 238 274699 272
rect 274389 210 274437 238
rect 274465 210 274499 238
rect 274527 210 274561 238
rect 274589 210 274623 238
rect 274651 210 274699 238
rect 274389 162 274699 210
rect 281529 299190 281839 299718
rect 281529 299162 281577 299190
rect 281605 299162 281639 299190
rect 281667 299162 281701 299190
rect 281729 299162 281763 299190
rect 281791 299162 281839 299190
rect 281529 299128 281839 299162
rect 281529 299100 281577 299128
rect 281605 299100 281639 299128
rect 281667 299100 281701 299128
rect 281729 299100 281763 299128
rect 281791 299100 281839 299128
rect 281529 299066 281839 299100
rect 281529 299038 281577 299066
rect 281605 299038 281639 299066
rect 281667 299038 281701 299066
rect 281729 299038 281763 299066
rect 281791 299038 281839 299066
rect 281529 299004 281839 299038
rect 281529 298976 281577 299004
rect 281605 298976 281639 299004
rect 281667 298976 281701 299004
rect 281729 298976 281763 299004
rect 281791 298976 281839 299004
rect 281529 290959 281839 298976
rect 281529 290931 281577 290959
rect 281605 290931 281639 290959
rect 281667 290931 281701 290959
rect 281729 290931 281763 290959
rect 281791 290931 281839 290959
rect 281529 290897 281839 290931
rect 281529 290869 281577 290897
rect 281605 290869 281639 290897
rect 281667 290869 281701 290897
rect 281729 290869 281763 290897
rect 281791 290869 281839 290897
rect 281529 290835 281839 290869
rect 281529 290807 281577 290835
rect 281605 290807 281639 290835
rect 281667 290807 281701 290835
rect 281729 290807 281763 290835
rect 281791 290807 281839 290835
rect 281529 290773 281839 290807
rect 281529 290745 281577 290773
rect 281605 290745 281639 290773
rect 281667 290745 281701 290773
rect 281729 290745 281763 290773
rect 281791 290745 281839 290773
rect 281529 281959 281839 290745
rect 281529 281931 281577 281959
rect 281605 281931 281639 281959
rect 281667 281931 281701 281959
rect 281729 281931 281763 281959
rect 281791 281931 281839 281959
rect 281529 281897 281839 281931
rect 281529 281869 281577 281897
rect 281605 281869 281639 281897
rect 281667 281869 281701 281897
rect 281729 281869 281763 281897
rect 281791 281869 281839 281897
rect 281529 281835 281839 281869
rect 281529 281807 281577 281835
rect 281605 281807 281639 281835
rect 281667 281807 281701 281835
rect 281729 281807 281763 281835
rect 281791 281807 281839 281835
rect 281529 281773 281839 281807
rect 281529 281745 281577 281773
rect 281605 281745 281639 281773
rect 281667 281745 281701 281773
rect 281729 281745 281763 281773
rect 281791 281745 281839 281773
rect 281529 272959 281839 281745
rect 281529 272931 281577 272959
rect 281605 272931 281639 272959
rect 281667 272931 281701 272959
rect 281729 272931 281763 272959
rect 281791 272931 281839 272959
rect 281529 272897 281839 272931
rect 281529 272869 281577 272897
rect 281605 272869 281639 272897
rect 281667 272869 281701 272897
rect 281729 272869 281763 272897
rect 281791 272869 281839 272897
rect 281529 272835 281839 272869
rect 281529 272807 281577 272835
rect 281605 272807 281639 272835
rect 281667 272807 281701 272835
rect 281729 272807 281763 272835
rect 281791 272807 281839 272835
rect 281529 272773 281839 272807
rect 281529 272745 281577 272773
rect 281605 272745 281639 272773
rect 281667 272745 281701 272773
rect 281729 272745 281763 272773
rect 281791 272745 281839 272773
rect 281529 263959 281839 272745
rect 281529 263931 281577 263959
rect 281605 263931 281639 263959
rect 281667 263931 281701 263959
rect 281729 263931 281763 263959
rect 281791 263931 281839 263959
rect 281529 263897 281839 263931
rect 281529 263869 281577 263897
rect 281605 263869 281639 263897
rect 281667 263869 281701 263897
rect 281729 263869 281763 263897
rect 281791 263869 281839 263897
rect 281529 263835 281839 263869
rect 281529 263807 281577 263835
rect 281605 263807 281639 263835
rect 281667 263807 281701 263835
rect 281729 263807 281763 263835
rect 281791 263807 281839 263835
rect 281529 263773 281839 263807
rect 281529 263745 281577 263773
rect 281605 263745 281639 263773
rect 281667 263745 281701 263773
rect 281729 263745 281763 263773
rect 281791 263745 281839 263773
rect 281529 254959 281839 263745
rect 281529 254931 281577 254959
rect 281605 254931 281639 254959
rect 281667 254931 281701 254959
rect 281729 254931 281763 254959
rect 281791 254931 281839 254959
rect 281529 254897 281839 254931
rect 281529 254869 281577 254897
rect 281605 254869 281639 254897
rect 281667 254869 281701 254897
rect 281729 254869 281763 254897
rect 281791 254869 281839 254897
rect 281529 254835 281839 254869
rect 281529 254807 281577 254835
rect 281605 254807 281639 254835
rect 281667 254807 281701 254835
rect 281729 254807 281763 254835
rect 281791 254807 281839 254835
rect 281529 254773 281839 254807
rect 281529 254745 281577 254773
rect 281605 254745 281639 254773
rect 281667 254745 281701 254773
rect 281729 254745 281763 254773
rect 281791 254745 281839 254773
rect 281529 245959 281839 254745
rect 281529 245931 281577 245959
rect 281605 245931 281639 245959
rect 281667 245931 281701 245959
rect 281729 245931 281763 245959
rect 281791 245931 281839 245959
rect 281529 245897 281839 245931
rect 281529 245869 281577 245897
rect 281605 245869 281639 245897
rect 281667 245869 281701 245897
rect 281729 245869 281763 245897
rect 281791 245869 281839 245897
rect 281529 245835 281839 245869
rect 281529 245807 281577 245835
rect 281605 245807 281639 245835
rect 281667 245807 281701 245835
rect 281729 245807 281763 245835
rect 281791 245807 281839 245835
rect 281529 245773 281839 245807
rect 281529 245745 281577 245773
rect 281605 245745 281639 245773
rect 281667 245745 281701 245773
rect 281729 245745 281763 245773
rect 281791 245745 281839 245773
rect 281529 236959 281839 245745
rect 281529 236931 281577 236959
rect 281605 236931 281639 236959
rect 281667 236931 281701 236959
rect 281729 236931 281763 236959
rect 281791 236931 281839 236959
rect 281529 236897 281839 236931
rect 281529 236869 281577 236897
rect 281605 236869 281639 236897
rect 281667 236869 281701 236897
rect 281729 236869 281763 236897
rect 281791 236869 281839 236897
rect 281529 236835 281839 236869
rect 281529 236807 281577 236835
rect 281605 236807 281639 236835
rect 281667 236807 281701 236835
rect 281729 236807 281763 236835
rect 281791 236807 281839 236835
rect 281529 236773 281839 236807
rect 281529 236745 281577 236773
rect 281605 236745 281639 236773
rect 281667 236745 281701 236773
rect 281729 236745 281763 236773
rect 281791 236745 281839 236773
rect 281529 227959 281839 236745
rect 281529 227931 281577 227959
rect 281605 227931 281639 227959
rect 281667 227931 281701 227959
rect 281729 227931 281763 227959
rect 281791 227931 281839 227959
rect 281529 227897 281839 227931
rect 281529 227869 281577 227897
rect 281605 227869 281639 227897
rect 281667 227869 281701 227897
rect 281729 227869 281763 227897
rect 281791 227869 281839 227897
rect 281529 227835 281839 227869
rect 281529 227807 281577 227835
rect 281605 227807 281639 227835
rect 281667 227807 281701 227835
rect 281729 227807 281763 227835
rect 281791 227807 281839 227835
rect 281529 227773 281839 227807
rect 281529 227745 281577 227773
rect 281605 227745 281639 227773
rect 281667 227745 281701 227773
rect 281729 227745 281763 227773
rect 281791 227745 281839 227773
rect 281529 218959 281839 227745
rect 281529 218931 281577 218959
rect 281605 218931 281639 218959
rect 281667 218931 281701 218959
rect 281729 218931 281763 218959
rect 281791 218931 281839 218959
rect 281529 218897 281839 218931
rect 281529 218869 281577 218897
rect 281605 218869 281639 218897
rect 281667 218869 281701 218897
rect 281729 218869 281763 218897
rect 281791 218869 281839 218897
rect 281529 218835 281839 218869
rect 281529 218807 281577 218835
rect 281605 218807 281639 218835
rect 281667 218807 281701 218835
rect 281729 218807 281763 218835
rect 281791 218807 281839 218835
rect 281529 218773 281839 218807
rect 281529 218745 281577 218773
rect 281605 218745 281639 218773
rect 281667 218745 281701 218773
rect 281729 218745 281763 218773
rect 281791 218745 281839 218773
rect 281529 209959 281839 218745
rect 281529 209931 281577 209959
rect 281605 209931 281639 209959
rect 281667 209931 281701 209959
rect 281729 209931 281763 209959
rect 281791 209931 281839 209959
rect 281529 209897 281839 209931
rect 281529 209869 281577 209897
rect 281605 209869 281639 209897
rect 281667 209869 281701 209897
rect 281729 209869 281763 209897
rect 281791 209869 281839 209897
rect 281529 209835 281839 209869
rect 281529 209807 281577 209835
rect 281605 209807 281639 209835
rect 281667 209807 281701 209835
rect 281729 209807 281763 209835
rect 281791 209807 281839 209835
rect 281529 209773 281839 209807
rect 281529 209745 281577 209773
rect 281605 209745 281639 209773
rect 281667 209745 281701 209773
rect 281729 209745 281763 209773
rect 281791 209745 281839 209773
rect 281529 200959 281839 209745
rect 281529 200931 281577 200959
rect 281605 200931 281639 200959
rect 281667 200931 281701 200959
rect 281729 200931 281763 200959
rect 281791 200931 281839 200959
rect 281529 200897 281839 200931
rect 281529 200869 281577 200897
rect 281605 200869 281639 200897
rect 281667 200869 281701 200897
rect 281729 200869 281763 200897
rect 281791 200869 281839 200897
rect 281529 200835 281839 200869
rect 281529 200807 281577 200835
rect 281605 200807 281639 200835
rect 281667 200807 281701 200835
rect 281729 200807 281763 200835
rect 281791 200807 281839 200835
rect 281529 200773 281839 200807
rect 281529 200745 281577 200773
rect 281605 200745 281639 200773
rect 281667 200745 281701 200773
rect 281729 200745 281763 200773
rect 281791 200745 281839 200773
rect 281529 191959 281839 200745
rect 281529 191931 281577 191959
rect 281605 191931 281639 191959
rect 281667 191931 281701 191959
rect 281729 191931 281763 191959
rect 281791 191931 281839 191959
rect 281529 191897 281839 191931
rect 281529 191869 281577 191897
rect 281605 191869 281639 191897
rect 281667 191869 281701 191897
rect 281729 191869 281763 191897
rect 281791 191869 281839 191897
rect 281529 191835 281839 191869
rect 281529 191807 281577 191835
rect 281605 191807 281639 191835
rect 281667 191807 281701 191835
rect 281729 191807 281763 191835
rect 281791 191807 281839 191835
rect 281529 191773 281839 191807
rect 281529 191745 281577 191773
rect 281605 191745 281639 191773
rect 281667 191745 281701 191773
rect 281729 191745 281763 191773
rect 281791 191745 281839 191773
rect 281529 182959 281839 191745
rect 281529 182931 281577 182959
rect 281605 182931 281639 182959
rect 281667 182931 281701 182959
rect 281729 182931 281763 182959
rect 281791 182931 281839 182959
rect 281529 182897 281839 182931
rect 281529 182869 281577 182897
rect 281605 182869 281639 182897
rect 281667 182869 281701 182897
rect 281729 182869 281763 182897
rect 281791 182869 281839 182897
rect 281529 182835 281839 182869
rect 281529 182807 281577 182835
rect 281605 182807 281639 182835
rect 281667 182807 281701 182835
rect 281729 182807 281763 182835
rect 281791 182807 281839 182835
rect 281529 182773 281839 182807
rect 281529 182745 281577 182773
rect 281605 182745 281639 182773
rect 281667 182745 281701 182773
rect 281729 182745 281763 182773
rect 281791 182745 281839 182773
rect 281529 173959 281839 182745
rect 281529 173931 281577 173959
rect 281605 173931 281639 173959
rect 281667 173931 281701 173959
rect 281729 173931 281763 173959
rect 281791 173931 281839 173959
rect 281529 173897 281839 173931
rect 281529 173869 281577 173897
rect 281605 173869 281639 173897
rect 281667 173869 281701 173897
rect 281729 173869 281763 173897
rect 281791 173869 281839 173897
rect 281529 173835 281839 173869
rect 281529 173807 281577 173835
rect 281605 173807 281639 173835
rect 281667 173807 281701 173835
rect 281729 173807 281763 173835
rect 281791 173807 281839 173835
rect 281529 173773 281839 173807
rect 281529 173745 281577 173773
rect 281605 173745 281639 173773
rect 281667 173745 281701 173773
rect 281729 173745 281763 173773
rect 281791 173745 281839 173773
rect 281529 164959 281839 173745
rect 281529 164931 281577 164959
rect 281605 164931 281639 164959
rect 281667 164931 281701 164959
rect 281729 164931 281763 164959
rect 281791 164931 281839 164959
rect 281529 164897 281839 164931
rect 281529 164869 281577 164897
rect 281605 164869 281639 164897
rect 281667 164869 281701 164897
rect 281729 164869 281763 164897
rect 281791 164869 281839 164897
rect 281529 164835 281839 164869
rect 281529 164807 281577 164835
rect 281605 164807 281639 164835
rect 281667 164807 281701 164835
rect 281729 164807 281763 164835
rect 281791 164807 281839 164835
rect 281529 164773 281839 164807
rect 281529 164745 281577 164773
rect 281605 164745 281639 164773
rect 281667 164745 281701 164773
rect 281729 164745 281763 164773
rect 281791 164745 281839 164773
rect 281529 155959 281839 164745
rect 281529 155931 281577 155959
rect 281605 155931 281639 155959
rect 281667 155931 281701 155959
rect 281729 155931 281763 155959
rect 281791 155931 281839 155959
rect 281529 155897 281839 155931
rect 281529 155869 281577 155897
rect 281605 155869 281639 155897
rect 281667 155869 281701 155897
rect 281729 155869 281763 155897
rect 281791 155869 281839 155897
rect 281529 155835 281839 155869
rect 281529 155807 281577 155835
rect 281605 155807 281639 155835
rect 281667 155807 281701 155835
rect 281729 155807 281763 155835
rect 281791 155807 281839 155835
rect 281529 155773 281839 155807
rect 281529 155745 281577 155773
rect 281605 155745 281639 155773
rect 281667 155745 281701 155773
rect 281729 155745 281763 155773
rect 281791 155745 281839 155773
rect 281529 146959 281839 155745
rect 281529 146931 281577 146959
rect 281605 146931 281639 146959
rect 281667 146931 281701 146959
rect 281729 146931 281763 146959
rect 281791 146931 281839 146959
rect 281529 146897 281839 146931
rect 281529 146869 281577 146897
rect 281605 146869 281639 146897
rect 281667 146869 281701 146897
rect 281729 146869 281763 146897
rect 281791 146869 281839 146897
rect 281529 146835 281839 146869
rect 281529 146807 281577 146835
rect 281605 146807 281639 146835
rect 281667 146807 281701 146835
rect 281729 146807 281763 146835
rect 281791 146807 281839 146835
rect 281529 146773 281839 146807
rect 281529 146745 281577 146773
rect 281605 146745 281639 146773
rect 281667 146745 281701 146773
rect 281729 146745 281763 146773
rect 281791 146745 281839 146773
rect 281529 137959 281839 146745
rect 281529 137931 281577 137959
rect 281605 137931 281639 137959
rect 281667 137931 281701 137959
rect 281729 137931 281763 137959
rect 281791 137931 281839 137959
rect 281529 137897 281839 137931
rect 281529 137869 281577 137897
rect 281605 137869 281639 137897
rect 281667 137869 281701 137897
rect 281729 137869 281763 137897
rect 281791 137869 281839 137897
rect 281529 137835 281839 137869
rect 281529 137807 281577 137835
rect 281605 137807 281639 137835
rect 281667 137807 281701 137835
rect 281729 137807 281763 137835
rect 281791 137807 281839 137835
rect 281529 137773 281839 137807
rect 281529 137745 281577 137773
rect 281605 137745 281639 137773
rect 281667 137745 281701 137773
rect 281729 137745 281763 137773
rect 281791 137745 281839 137773
rect 281529 128959 281839 137745
rect 281529 128931 281577 128959
rect 281605 128931 281639 128959
rect 281667 128931 281701 128959
rect 281729 128931 281763 128959
rect 281791 128931 281839 128959
rect 281529 128897 281839 128931
rect 281529 128869 281577 128897
rect 281605 128869 281639 128897
rect 281667 128869 281701 128897
rect 281729 128869 281763 128897
rect 281791 128869 281839 128897
rect 281529 128835 281839 128869
rect 281529 128807 281577 128835
rect 281605 128807 281639 128835
rect 281667 128807 281701 128835
rect 281729 128807 281763 128835
rect 281791 128807 281839 128835
rect 281529 128773 281839 128807
rect 281529 128745 281577 128773
rect 281605 128745 281639 128773
rect 281667 128745 281701 128773
rect 281729 128745 281763 128773
rect 281791 128745 281839 128773
rect 281529 119959 281839 128745
rect 281529 119931 281577 119959
rect 281605 119931 281639 119959
rect 281667 119931 281701 119959
rect 281729 119931 281763 119959
rect 281791 119931 281839 119959
rect 281529 119897 281839 119931
rect 281529 119869 281577 119897
rect 281605 119869 281639 119897
rect 281667 119869 281701 119897
rect 281729 119869 281763 119897
rect 281791 119869 281839 119897
rect 281529 119835 281839 119869
rect 281529 119807 281577 119835
rect 281605 119807 281639 119835
rect 281667 119807 281701 119835
rect 281729 119807 281763 119835
rect 281791 119807 281839 119835
rect 281529 119773 281839 119807
rect 281529 119745 281577 119773
rect 281605 119745 281639 119773
rect 281667 119745 281701 119773
rect 281729 119745 281763 119773
rect 281791 119745 281839 119773
rect 281529 110959 281839 119745
rect 281529 110931 281577 110959
rect 281605 110931 281639 110959
rect 281667 110931 281701 110959
rect 281729 110931 281763 110959
rect 281791 110931 281839 110959
rect 281529 110897 281839 110931
rect 281529 110869 281577 110897
rect 281605 110869 281639 110897
rect 281667 110869 281701 110897
rect 281729 110869 281763 110897
rect 281791 110869 281839 110897
rect 281529 110835 281839 110869
rect 281529 110807 281577 110835
rect 281605 110807 281639 110835
rect 281667 110807 281701 110835
rect 281729 110807 281763 110835
rect 281791 110807 281839 110835
rect 281529 110773 281839 110807
rect 281529 110745 281577 110773
rect 281605 110745 281639 110773
rect 281667 110745 281701 110773
rect 281729 110745 281763 110773
rect 281791 110745 281839 110773
rect 281529 101959 281839 110745
rect 281529 101931 281577 101959
rect 281605 101931 281639 101959
rect 281667 101931 281701 101959
rect 281729 101931 281763 101959
rect 281791 101931 281839 101959
rect 281529 101897 281839 101931
rect 281529 101869 281577 101897
rect 281605 101869 281639 101897
rect 281667 101869 281701 101897
rect 281729 101869 281763 101897
rect 281791 101869 281839 101897
rect 281529 101835 281839 101869
rect 281529 101807 281577 101835
rect 281605 101807 281639 101835
rect 281667 101807 281701 101835
rect 281729 101807 281763 101835
rect 281791 101807 281839 101835
rect 281529 101773 281839 101807
rect 281529 101745 281577 101773
rect 281605 101745 281639 101773
rect 281667 101745 281701 101773
rect 281729 101745 281763 101773
rect 281791 101745 281839 101773
rect 281529 92959 281839 101745
rect 281529 92931 281577 92959
rect 281605 92931 281639 92959
rect 281667 92931 281701 92959
rect 281729 92931 281763 92959
rect 281791 92931 281839 92959
rect 281529 92897 281839 92931
rect 281529 92869 281577 92897
rect 281605 92869 281639 92897
rect 281667 92869 281701 92897
rect 281729 92869 281763 92897
rect 281791 92869 281839 92897
rect 281529 92835 281839 92869
rect 281529 92807 281577 92835
rect 281605 92807 281639 92835
rect 281667 92807 281701 92835
rect 281729 92807 281763 92835
rect 281791 92807 281839 92835
rect 281529 92773 281839 92807
rect 281529 92745 281577 92773
rect 281605 92745 281639 92773
rect 281667 92745 281701 92773
rect 281729 92745 281763 92773
rect 281791 92745 281839 92773
rect 281529 83959 281839 92745
rect 281529 83931 281577 83959
rect 281605 83931 281639 83959
rect 281667 83931 281701 83959
rect 281729 83931 281763 83959
rect 281791 83931 281839 83959
rect 281529 83897 281839 83931
rect 281529 83869 281577 83897
rect 281605 83869 281639 83897
rect 281667 83869 281701 83897
rect 281729 83869 281763 83897
rect 281791 83869 281839 83897
rect 281529 83835 281839 83869
rect 281529 83807 281577 83835
rect 281605 83807 281639 83835
rect 281667 83807 281701 83835
rect 281729 83807 281763 83835
rect 281791 83807 281839 83835
rect 281529 83773 281839 83807
rect 281529 83745 281577 83773
rect 281605 83745 281639 83773
rect 281667 83745 281701 83773
rect 281729 83745 281763 83773
rect 281791 83745 281839 83773
rect 281529 74959 281839 83745
rect 281529 74931 281577 74959
rect 281605 74931 281639 74959
rect 281667 74931 281701 74959
rect 281729 74931 281763 74959
rect 281791 74931 281839 74959
rect 281529 74897 281839 74931
rect 281529 74869 281577 74897
rect 281605 74869 281639 74897
rect 281667 74869 281701 74897
rect 281729 74869 281763 74897
rect 281791 74869 281839 74897
rect 281529 74835 281839 74869
rect 281529 74807 281577 74835
rect 281605 74807 281639 74835
rect 281667 74807 281701 74835
rect 281729 74807 281763 74835
rect 281791 74807 281839 74835
rect 281529 74773 281839 74807
rect 281529 74745 281577 74773
rect 281605 74745 281639 74773
rect 281667 74745 281701 74773
rect 281729 74745 281763 74773
rect 281791 74745 281839 74773
rect 281529 65959 281839 74745
rect 281529 65931 281577 65959
rect 281605 65931 281639 65959
rect 281667 65931 281701 65959
rect 281729 65931 281763 65959
rect 281791 65931 281839 65959
rect 281529 65897 281839 65931
rect 281529 65869 281577 65897
rect 281605 65869 281639 65897
rect 281667 65869 281701 65897
rect 281729 65869 281763 65897
rect 281791 65869 281839 65897
rect 281529 65835 281839 65869
rect 281529 65807 281577 65835
rect 281605 65807 281639 65835
rect 281667 65807 281701 65835
rect 281729 65807 281763 65835
rect 281791 65807 281839 65835
rect 281529 65773 281839 65807
rect 281529 65745 281577 65773
rect 281605 65745 281639 65773
rect 281667 65745 281701 65773
rect 281729 65745 281763 65773
rect 281791 65745 281839 65773
rect 281529 56959 281839 65745
rect 281529 56931 281577 56959
rect 281605 56931 281639 56959
rect 281667 56931 281701 56959
rect 281729 56931 281763 56959
rect 281791 56931 281839 56959
rect 281529 56897 281839 56931
rect 281529 56869 281577 56897
rect 281605 56869 281639 56897
rect 281667 56869 281701 56897
rect 281729 56869 281763 56897
rect 281791 56869 281839 56897
rect 281529 56835 281839 56869
rect 281529 56807 281577 56835
rect 281605 56807 281639 56835
rect 281667 56807 281701 56835
rect 281729 56807 281763 56835
rect 281791 56807 281839 56835
rect 281529 56773 281839 56807
rect 281529 56745 281577 56773
rect 281605 56745 281639 56773
rect 281667 56745 281701 56773
rect 281729 56745 281763 56773
rect 281791 56745 281839 56773
rect 281529 47959 281839 56745
rect 281529 47931 281577 47959
rect 281605 47931 281639 47959
rect 281667 47931 281701 47959
rect 281729 47931 281763 47959
rect 281791 47931 281839 47959
rect 281529 47897 281839 47931
rect 281529 47869 281577 47897
rect 281605 47869 281639 47897
rect 281667 47869 281701 47897
rect 281729 47869 281763 47897
rect 281791 47869 281839 47897
rect 281529 47835 281839 47869
rect 281529 47807 281577 47835
rect 281605 47807 281639 47835
rect 281667 47807 281701 47835
rect 281729 47807 281763 47835
rect 281791 47807 281839 47835
rect 281529 47773 281839 47807
rect 281529 47745 281577 47773
rect 281605 47745 281639 47773
rect 281667 47745 281701 47773
rect 281729 47745 281763 47773
rect 281791 47745 281839 47773
rect 281529 38959 281839 47745
rect 281529 38931 281577 38959
rect 281605 38931 281639 38959
rect 281667 38931 281701 38959
rect 281729 38931 281763 38959
rect 281791 38931 281839 38959
rect 281529 38897 281839 38931
rect 281529 38869 281577 38897
rect 281605 38869 281639 38897
rect 281667 38869 281701 38897
rect 281729 38869 281763 38897
rect 281791 38869 281839 38897
rect 281529 38835 281839 38869
rect 281529 38807 281577 38835
rect 281605 38807 281639 38835
rect 281667 38807 281701 38835
rect 281729 38807 281763 38835
rect 281791 38807 281839 38835
rect 281529 38773 281839 38807
rect 281529 38745 281577 38773
rect 281605 38745 281639 38773
rect 281667 38745 281701 38773
rect 281729 38745 281763 38773
rect 281791 38745 281839 38773
rect 281529 29959 281839 38745
rect 281529 29931 281577 29959
rect 281605 29931 281639 29959
rect 281667 29931 281701 29959
rect 281729 29931 281763 29959
rect 281791 29931 281839 29959
rect 281529 29897 281839 29931
rect 281529 29869 281577 29897
rect 281605 29869 281639 29897
rect 281667 29869 281701 29897
rect 281729 29869 281763 29897
rect 281791 29869 281839 29897
rect 281529 29835 281839 29869
rect 281529 29807 281577 29835
rect 281605 29807 281639 29835
rect 281667 29807 281701 29835
rect 281729 29807 281763 29835
rect 281791 29807 281839 29835
rect 281529 29773 281839 29807
rect 281529 29745 281577 29773
rect 281605 29745 281639 29773
rect 281667 29745 281701 29773
rect 281729 29745 281763 29773
rect 281791 29745 281839 29773
rect 281529 20959 281839 29745
rect 281529 20931 281577 20959
rect 281605 20931 281639 20959
rect 281667 20931 281701 20959
rect 281729 20931 281763 20959
rect 281791 20931 281839 20959
rect 281529 20897 281839 20931
rect 281529 20869 281577 20897
rect 281605 20869 281639 20897
rect 281667 20869 281701 20897
rect 281729 20869 281763 20897
rect 281791 20869 281839 20897
rect 281529 20835 281839 20869
rect 281529 20807 281577 20835
rect 281605 20807 281639 20835
rect 281667 20807 281701 20835
rect 281729 20807 281763 20835
rect 281791 20807 281839 20835
rect 281529 20773 281839 20807
rect 281529 20745 281577 20773
rect 281605 20745 281639 20773
rect 281667 20745 281701 20773
rect 281729 20745 281763 20773
rect 281791 20745 281839 20773
rect 281529 11959 281839 20745
rect 281529 11931 281577 11959
rect 281605 11931 281639 11959
rect 281667 11931 281701 11959
rect 281729 11931 281763 11959
rect 281791 11931 281839 11959
rect 281529 11897 281839 11931
rect 281529 11869 281577 11897
rect 281605 11869 281639 11897
rect 281667 11869 281701 11897
rect 281729 11869 281763 11897
rect 281791 11869 281839 11897
rect 281529 11835 281839 11869
rect 281529 11807 281577 11835
rect 281605 11807 281639 11835
rect 281667 11807 281701 11835
rect 281729 11807 281763 11835
rect 281791 11807 281839 11835
rect 281529 11773 281839 11807
rect 281529 11745 281577 11773
rect 281605 11745 281639 11773
rect 281667 11745 281701 11773
rect 281729 11745 281763 11773
rect 281791 11745 281839 11773
rect 281529 2959 281839 11745
rect 281529 2931 281577 2959
rect 281605 2931 281639 2959
rect 281667 2931 281701 2959
rect 281729 2931 281763 2959
rect 281791 2931 281839 2959
rect 281529 2897 281839 2931
rect 281529 2869 281577 2897
rect 281605 2869 281639 2897
rect 281667 2869 281701 2897
rect 281729 2869 281763 2897
rect 281791 2869 281839 2897
rect 281529 2835 281839 2869
rect 281529 2807 281577 2835
rect 281605 2807 281639 2835
rect 281667 2807 281701 2835
rect 281729 2807 281763 2835
rect 281791 2807 281839 2835
rect 281529 2773 281839 2807
rect 281529 2745 281577 2773
rect 281605 2745 281639 2773
rect 281667 2745 281701 2773
rect 281729 2745 281763 2773
rect 281791 2745 281839 2773
rect 281529 904 281839 2745
rect 281529 876 281577 904
rect 281605 876 281639 904
rect 281667 876 281701 904
rect 281729 876 281763 904
rect 281791 876 281839 904
rect 281529 842 281839 876
rect 281529 814 281577 842
rect 281605 814 281639 842
rect 281667 814 281701 842
rect 281729 814 281763 842
rect 281791 814 281839 842
rect 281529 780 281839 814
rect 281529 752 281577 780
rect 281605 752 281639 780
rect 281667 752 281701 780
rect 281729 752 281763 780
rect 281791 752 281839 780
rect 281529 718 281839 752
rect 281529 690 281577 718
rect 281605 690 281639 718
rect 281667 690 281701 718
rect 281729 690 281763 718
rect 281791 690 281839 718
rect 281529 162 281839 690
rect 283389 299670 283699 299718
rect 283389 299642 283437 299670
rect 283465 299642 283499 299670
rect 283527 299642 283561 299670
rect 283589 299642 283623 299670
rect 283651 299642 283699 299670
rect 283389 299608 283699 299642
rect 283389 299580 283437 299608
rect 283465 299580 283499 299608
rect 283527 299580 283561 299608
rect 283589 299580 283623 299608
rect 283651 299580 283699 299608
rect 283389 299546 283699 299580
rect 283389 299518 283437 299546
rect 283465 299518 283499 299546
rect 283527 299518 283561 299546
rect 283589 299518 283623 299546
rect 283651 299518 283699 299546
rect 283389 299484 283699 299518
rect 283389 299456 283437 299484
rect 283465 299456 283499 299484
rect 283527 299456 283561 299484
rect 283589 299456 283623 299484
rect 283651 299456 283699 299484
rect 283389 293959 283699 299456
rect 283389 293931 283437 293959
rect 283465 293931 283499 293959
rect 283527 293931 283561 293959
rect 283589 293931 283623 293959
rect 283651 293931 283699 293959
rect 283389 293897 283699 293931
rect 283389 293869 283437 293897
rect 283465 293869 283499 293897
rect 283527 293869 283561 293897
rect 283589 293869 283623 293897
rect 283651 293869 283699 293897
rect 283389 293835 283699 293869
rect 283389 293807 283437 293835
rect 283465 293807 283499 293835
rect 283527 293807 283561 293835
rect 283589 293807 283623 293835
rect 283651 293807 283699 293835
rect 283389 293773 283699 293807
rect 283389 293745 283437 293773
rect 283465 293745 283499 293773
rect 283527 293745 283561 293773
rect 283589 293745 283623 293773
rect 283651 293745 283699 293773
rect 283389 284959 283699 293745
rect 283389 284931 283437 284959
rect 283465 284931 283499 284959
rect 283527 284931 283561 284959
rect 283589 284931 283623 284959
rect 283651 284931 283699 284959
rect 283389 284897 283699 284931
rect 283389 284869 283437 284897
rect 283465 284869 283499 284897
rect 283527 284869 283561 284897
rect 283589 284869 283623 284897
rect 283651 284869 283699 284897
rect 283389 284835 283699 284869
rect 283389 284807 283437 284835
rect 283465 284807 283499 284835
rect 283527 284807 283561 284835
rect 283589 284807 283623 284835
rect 283651 284807 283699 284835
rect 283389 284773 283699 284807
rect 283389 284745 283437 284773
rect 283465 284745 283499 284773
rect 283527 284745 283561 284773
rect 283589 284745 283623 284773
rect 283651 284745 283699 284773
rect 283389 275959 283699 284745
rect 283389 275931 283437 275959
rect 283465 275931 283499 275959
rect 283527 275931 283561 275959
rect 283589 275931 283623 275959
rect 283651 275931 283699 275959
rect 283389 275897 283699 275931
rect 283389 275869 283437 275897
rect 283465 275869 283499 275897
rect 283527 275869 283561 275897
rect 283589 275869 283623 275897
rect 283651 275869 283699 275897
rect 283389 275835 283699 275869
rect 283389 275807 283437 275835
rect 283465 275807 283499 275835
rect 283527 275807 283561 275835
rect 283589 275807 283623 275835
rect 283651 275807 283699 275835
rect 283389 275773 283699 275807
rect 283389 275745 283437 275773
rect 283465 275745 283499 275773
rect 283527 275745 283561 275773
rect 283589 275745 283623 275773
rect 283651 275745 283699 275773
rect 283389 266959 283699 275745
rect 283389 266931 283437 266959
rect 283465 266931 283499 266959
rect 283527 266931 283561 266959
rect 283589 266931 283623 266959
rect 283651 266931 283699 266959
rect 283389 266897 283699 266931
rect 283389 266869 283437 266897
rect 283465 266869 283499 266897
rect 283527 266869 283561 266897
rect 283589 266869 283623 266897
rect 283651 266869 283699 266897
rect 283389 266835 283699 266869
rect 283389 266807 283437 266835
rect 283465 266807 283499 266835
rect 283527 266807 283561 266835
rect 283589 266807 283623 266835
rect 283651 266807 283699 266835
rect 283389 266773 283699 266807
rect 283389 266745 283437 266773
rect 283465 266745 283499 266773
rect 283527 266745 283561 266773
rect 283589 266745 283623 266773
rect 283651 266745 283699 266773
rect 283389 257959 283699 266745
rect 283389 257931 283437 257959
rect 283465 257931 283499 257959
rect 283527 257931 283561 257959
rect 283589 257931 283623 257959
rect 283651 257931 283699 257959
rect 283389 257897 283699 257931
rect 283389 257869 283437 257897
rect 283465 257869 283499 257897
rect 283527 257869 283561 257897
rect 283589 257869 283623 257897
rect 283651 257869 283699 257897
rect 283389 257835 283699 257869
rect 283389 257807 283437 257835
rect 283465 257807 283499 257835
rect 283527 257807 283561 257835
rect 283589 257807 283623 257835
rect 283651 257807 283699 257835
rect 283389 257773 283699 257807
rect 283389 257745 283437 257773
rect 283465 257745 283499 257773
rect 283527 257745 283561 257773
rect 283589 257745 283623 257773
rect 283651 257745 283699 257773
rect 283389 248959 283699 257745
rect 283389 248931 283437 248959
rect 283465 248931 283499 248959
rect 283527 248931 283561 248959
rect 283589 248931 283623 248959
rect 283651 248931 283699 248959
rect 283389 248897 283699 248931
rect 283389 248869 283437 248897
rect 283465 248869 283499 248897
rect 283527 248869 283561 248897
rect 283589 248869 283623 248897
rect 283651 248869 283699 248897
rect 283389 248835 283699 248869
rect 283389 248807 283437 248835
rect 283465 248807 283499 248835
rect 283527 248807 283561 248835
rect 283589 248807 283623 248835
rect 283651 248807 283699 248835
rect 283389 248773 283699 248807
rect 283389 248745 283437 248773
rect 283465 248745 283499 248773
rect 283527 248745 283561 248773
rect 283589 248745 283623 248773
rect 283651 248745 283699 248773
rect 283389 239959 283699 248745
rect 283389 239931 283437 239959
rect 283465 239931 283499 239959
rect 283527 239931 283561 239959
rect 283589 239931 283623 239959
rect 283651 239931 283699 239959
rect 283389 239897 283699 239931
rect 283389 239869 283437 239897
rect 283465 239869 283499 239897
rect 283527 239869 283561 239897
rect 283589 239869 283623 239897
rect 283651 239869 283699 239897
rect 283389 239835 283699 239869
rect 283389 239807 283437 239835
rect 283465 239807 283499 239835
rect 283527 239807 283561 239835
rect 283589 239807 283623 239835
rect 283651 239807 283699 239835
rect 283389 239773 283699 239807
rect 283389 239745 283437 239773
rect 283465 239745 283499 239773
rect 283527 239745 283561 239773
rect 283589 239745 283623 239773
rect 283651 239745 283699 239773
rect 283389 230959 283699 239745
rect 283389 230931 283437 230959
rect 283465 230931 283499 230959
rect 283527 230931 283561 230959
rect 283589 230931 283623 230959
rect 283651 230931 283699 230959
rect 283389 230897 283699 230931
rect 283389 230869 283437 230897
rect 283465 230869 283499 230897
rect 283527 230869 283561 230897
rect 283589 230869 283623 230897
rect 283651 230869 283699 230897
rect 283389 230835 283699 230869
rect 283389 230807 283437 230835
rect 283465 230807 283499 230835
rect 283527 230807 283561 230835
rect 283589 230807 283623 230835
rect 283651 230807 283699 230835
rect 283389 230773 283699 230807
rect 283389 230745 283437 230773
rect 283465 230745 283499 230773
rect 283527 230745 283561 230773
rect 283589 230745 283623 230773
rect 283651 230745 283699 230773
rect 283389 221959 283699 230745
rect 283389 221931 283437 221959
rect 283465 221931 283499 221959
rect 283527 221931 283561 221959
rect 283589 221931 283623 221959
rect 283651 221931 283699 221959
rect 283389 221897 283699 221931
rect 283389 221869 283437 221897
rect 283465 221869 283499 221897
rect 283527 221869 283561 221897
rect 283589 221869 283623 221897
rect 283651 221869 283699 221897
rect 283389 221835 283699 221869
rect 283389 221807 283437 221835
rect 283465 221807 283499 221835
rect 283527 221807 283561 221835
rect 283589 221807 283623 221835
rect 283651 221807 283699 221835
rect 283389 221773 283699 221807
rect 283389 221745 283437 221773
rect 283465 221745 283499 221773
rect 283527 221745 283561 221773
rect 283589 221745 283623 221773
rect 283651 221745 283699 221773
rect 283389 212959 283699 221745
rect 283389 212931 283437 212959
rect 283465 212931 283499 212959
rect 283527 212931 283561 212959
rect 283589 212931 283623 212959
rect 283651 212931 283699 212959
rect 283389 212897 283699 212931
rect 283389 212869 283437 212897
rect 283465 212869 283499 212897
rect 283527 212869 283561 212897
rect 283589 212869 283623 212897
rect 283651 212869 283699 212897
rect 283389 212835 283699 212869
rect 283389 212807 283437 212835
rect 283465 212807 283499 212835
rect 283527 212807 283561 212835
rect 283589 212807 283623 212835
rect 283651 212807 283699 212835
rect 283389 212773 283699 212807
rect 283389 212745 283437 212773
rect 283465 212745 283499 212773
rect 283527 212745 283561 212773
rect 283589 212745 283623 212773
rect 283651 212745 283699 212773
rect 283389 203959 283699 212745
rect 283389 203931 283437 203959
rect 283465 203931 283499 203959
rect 283527 203931 283561 203959
rect 283589 203931 283623 203959
rect 283651 203931 283699 203959
rect 283389 203897 283699 203931
rect 283389 203869 283437 203897
rect 283465 203869 283499 203897
rect 283527 203869 283561 203897
rect 283589 203869 283623 203897
rect 283651 203869 283699 203897
rect 283389 203835 283699 203869
rect 283389 203807 283437 203835
rect 283465 203807 283499 203835
rect 283527 203807 283561 203835
rect 283589 203807 283623 203835
rect 283651 203807 283699 203835
rect 283389 203773 283699 203807
rect 283389 203745 283437 203773
rect 283465 203745 283499 203773
rect 283527 203745 283561 203773
rect 283589 203745 283623 203773
rect 283651 203745 283699 203773
rect 283389 194959 283699 203745
rect 283389 194931 283437 194959
rect 283465 194931 283499 194959
rect 283527 194931 283561 194959
rect 283589 194931 283623 194959
rect 283651 194931 283699 194959
rect 283389 194897 283699 194931
rect 283389 194869 283437 194897
rect 283465 194869 283499 194897
rect 283527 194869 283561 194897
rect 283589 194869 283623 194897
rect 283651 194869 283699 194897
rect 283389 194835 283699 194869
rect 283389 194807 283437 194835
rect 283465 194807 283499 194835
rect 283527 194807 283561 194835
rect 283589 194807 283623 194835
rect 283651 194807 283699 194835
rect 283389 194773 283699 194807
rect 283389 194745 283437 194773
rect 283465 194745 283499 194773
rect 283527 194745 283561 194773
rect 283589 194745 283623 194773
rect 283651 194745 283699 194773
rect 283389 185959 283699 194745
rect 283389 185931 283437 185959
rect 283465 185931 283499 185959
rect 283527 185931 283561 185959
rect 283589 185931 283623 185959
rect 283651 185931 283699 185959
rect 283389 185897 283699 185931
rect 283389 185869 283437 185897
rect 283465 185869 283499 185897
rect 283527 185869 283561 185897
rect 283589 185869 283623 185897
rect 283651 185869 283699 185897
rect 283389 185835 283699 185869
rect 283389 185807 283437 185835
rect 283465 185807 283499 185835
rect 283527 185807 283561 185835
rect 283589 185807 283623 185835
rect 283651 185807 283699 185835
rect 283389 185773 283699 185807
rect 283389 185745 283437 185773
rect 283465 185745 283499 185773
rect 283527 185745 283561 185773
rect 283589 185745 283623 185773
rect 283651 185745 283699 185773
rect 283389 176959 283699 185745
rect 283389 176931 283437 176959
rect 283465 176931 283499 176959
rect 283527 176931 283561 176959
rect 283589 176931 283623 176959
rect 283651 176931 283699 176959
rect 283389 176897 283699 176931
rect 283389 176869 283437 176897
rect 283465 176869 283499 176897
rect 283527 176869 283561 176897
rect 283589 176869 283623 176897
rect 283651 176869 283699 176897
rect 283389 176835 283699 176869
rect 283389 176807 283437 176835
rect 283465 176807 283499 176835
rect 283527 176807 283561 176835
rect 283589 176807 283623 176835
rect 283651 176807 283699 176835
rect 283389 176773 283699 176807
rect 283389 176745 283437 176773
rect 283465 176745 283499 176773
rect 283527 176745 283561 176773
rect 283589 176745 283623 176773
rect 283651 176745 283699 176773
rect 283389 167959 283699 176745
rect 283389 167931 283437 167959
rect 283465 167931 283499 167959
rect 283527 167931 283561 167959
rect 283589 167931 283623 167959
rect 283651 167931 283699 167959
rect 283389 167897 283699 167931
rect 283389 167869 283437 167897
rect 283465 167869 283499 167897
rect 283527 167869 283561 167897
rect 283589 167869 283623 167897
rect 283651 167869 283699 167897
rect 283389 167835 283699 167869
rect 283389 167807 283437 167835
rect 283465 167807 283499 167835
rect 283527 167807 283561 167835
rect 283589 167807 283623 167835
rect 283651 167807 283699 167835
rect 283389 167773 283699 167807
rect 283389 167745 283437 167773
rect 283465 167745 283499 167773
rect 283527 167745 283561 167773
rect 283589 167745 283623 167773
rect 283651 167745 283699 167773
rect 283389 158959 283699 167745
rect 283389 158931 283437 158959
rect 283465 158931 283499 158959
rect 283527 158931 283561 158959
rect 283589 158931 283623 158959
rect 283651 158931 283699 158959
rect 283389 158897 283699 158931
rect 283389 158869 283437 158897
rect 283465 158869 283499 158897
rect 283527 158869 283561 158897
rect 283589 158869 283623 158897
rect 283651 158869 283699 158897
rect 283389 158835 283699 158869
rect 283389 158807 283437 158835
rect 283465 158807 283499 158835
rect 283527 158807 283561 158835
rect 283589 158807 283623 158835
rect 283651 158807 283699 158835
rect 283389 158773 283699 158807
rect 283389 158745 283437 158773
rect 283465 158745 283499 158773
rect 283527 158745 283561 158773
rect 283589 158745 283623 158773
rect 283651 158745 283699 158773
rect 283389 149959 283699 158745
rect 283389 149931 283437 149959
rect 283465 149931 283499 149959
rect 283527 149931 283561 149959
rect 283589 149931 283623 149959
rect 283651 149931 283699 149959
rect 283389 149897 283699 149931
rect 283389 149869 283437 149897
rect 283465 149869 283499 149897
rect 283527 149869 283561 149897
rect 283589 149869 283623 149897
rect 283651 149869 283699 149897
rect 283389 149835 283699 149869
rect 283389 149807 283437 149835
rect 283465 149807 283499 149835
rect 283527 149807 283561 149835
rect 283589 149807 283623 149835
rect 283651 149807 283699 149835
rect 283389 149773 283699 149807
rect 283389 149745 283437 149773
rect 283465 149745 283499 149773
rect 283527 149745 283561 149773
rect 283589 149745 283623 149773
rect 283651 149745 283699 149773
rect 283389 140959 283699 149745
rect 283389 140931 283437 140959
rect 283465 140931 283499 140959
rect 283527 140931 283561 140959
rect 283589 140931 283623 140959
rect 283651 140931 283699 140959
rect 283389 140897 283699 140931
rect 283389 140869 283437 140897
rect 283465 140869 283499 140897
rect 283527 140869 283561 140897
rect 283589 140869 283623 140897
rect 283651 140869 283699 140897
rect 283389 140835 283699 140869
rect 283389 140807 283437 140835
rect 283465 140807 283499 140835
rect 283527 140807 283561 140835
rect 283589 140807 283623 140835
rect 283651 140807 283699 140835
rect 283389 140773 283699 140807
rect 283389 140745 283437 140773
rect 283465 140745 283499 140773
rect 283527 140745 283561 140773
rect 283589 140745 283623 140773
rect 283651 140745 283699 140773
rect 283389 131959 283699 140745
rect 283389 131931 283437 131959
rect 283465 131931 283499 131959
rect 283527 131931 283561 131959
rect 283589 131931 283623 131959
rect 283651 131931 283699 131959
rect 283389 131897 283699 131931
rect 283389 131869 283437 131897
rect 283465 131869 283499 131897
rect 283527 131869 283561 131897
rect 283589 131869 283623 131897
rect 283651 131869 283699 131897
rect 283389 131835 283699 131869
rect 283389 131807 283437 131835
rect 283465 131807 283499 131835
rect 283527 131807 283561 131835
rect 283589 131807 283623 131835
rect 283651 131807 283699 131835
rect 283389 131773 283699 131807
rect 283389 131745 283437 131773
rect 283465 131745 283499 131773
rect 283527 131745 283561 131773
rect 283589 131745 283623 131773
rect 283651 131745 283699 131773
rect 283389 122959 283699 131745
rect 283389 122931 283437 122959
rect 283465 122931 283499 122959
rect 283527 122931 283561 122959
rect 283589 122931 283623 122959
rect 283651 122931 283699 122959
rect 283389 122897 283699 122931
rect 283389 122869 283437 122897
rect 283465 122869 283499 122897
rect 283527 122869 283561 122897
rect 283589 122869 283623 122897
rect 283651 122869 283699 122897
rect 283389 122835 283699 122869
rect 283389 122807 283437 122835
rect 283465 122807 283499 122835
rect 283527 122807 283561 122835
rect 283589 122807 283623 122835
rect 283651 122807 283699 122835
rect 283389 122773 283699 122807
rect 283389 122745 283437 122773
rect 283465 122745 283499 122773
rect 283527 122745 283561 122773
rect 283589 122745 283623 122773
rect 283651 122745 283699 122773
rect 283389 113959 283699 122745
rect 283389 113931 283437 113959
rect 283465 113931 283499 113959
rect 283527 113931 283561 113959
rect 283589 113931 283623 113959
rect 283651 113931 283699 113959
rect 283389 113897 283699 113931
rect 283389 113869 283437 113897
rect 283465 113869 283499 113897
rect 283527 113869 283561 113897
rect 283589 113869 283623 113897
rect 283651 113869 283699 113897
rect 283389 113835 283699 113869
rect 283389 113807 283437 113835
rect 283465 113807 283499 113835
rect 283527 113807 283561 113835
rect 283589 113807 283623 113835
rect 283651 113807 283699 113835
rect 283389 113773 283699 113807
rect 283389 113745 283437 113773
rect 283465 113745 283499 113773
rect 283527 113745 283561 113773
rect 283589 113745 283623 113773
rect 283651 113745 283699 113773
rect 283389 104959 283699 113745
rect 283389 104931 283437 104959
rect 283465 104931 283499 104959
rect 283527 104931 283561 104959
rect 283589 104931 283623 104959
rect 283651 104931 283699 104959
rect 283389 104897 283699 104931
rect 283389 104869 283437 104897
rect 283465 104869 283499 104897
rect 283527 104869 283561 104897
rect 283589 104869 283623 104897
rect 283651 104869 283699 104897
rect 283389 104835 283699 104869
rect 283389 104807 283437 104835
rect 283465 104807 283499 104835
rect 283527 104807 283561 104835
rect 283589 104807 283623 104835
rect 283651 104807 283699 104835
rect 283389 104773 283699 104807
rect 283389 104745 283437 104773
rect 283465 104745 283499 104773
rect 283527 104745 283561 104773
rect 283589 104745 283623 104773
rect 283651 104745 283699 104773
rect 283389 95959 283699 104745
rect 283389 95931 283437 95959
rect 283465 95931 283499 95959
rect 283527 95931 283561 95959
rect 283589 95931 283623 95959
rect 283651 95931 283699 95959
rect 283389 95897 283699 95931
rect 283389 95869 283437 95897
rect 283465 95869 283499 95897
rect 283527 95869 283561 95897
rect 283589 95869 283623 95897
rect 283651 95869 283699 95897
rect 283389 95835 283699 95869
rect 283389 95807 283437 95835
rect 283465 95807 283499 95835
rect 283527 95807 283561 95835
rect 283589 95807 283623 95835
rect 283651 95807 283699 95835
rect 283389 95773 283699 95807
rect 283389 95745 283437 95773
rect 283465 95745 283499 95773
rect 283527 95745 283561 95773
rect 283589 95745 283623 95773
rect 283651 95745 283699 95773
rect 283389 86959 283699 95745
rect 283389 86931 283437 86959
rect 283465 86931 283499 86959
rect 283527 86931 283561 86959
rect 283589 86931 283623 86959
rect 283651 86931 283699 86959
rect 283389 86897 283699 86931
rect 283389 86869 283437 86897
rect 283465 86869 283499 86897
rect 283527 86869 283561 86897
rect 283589 86869 283623 86897
rect 283651 86869 283699 86897
rect 283389 86835 283699 86869
rect 283389 86807 283437 86835
rect 283465 86807 283499 86835
rect 283527 86807 283561 86835
rect 283589 86807 283623 86835
rect 283651 86807 283699 86835
rect 283389 86773 283699 86807
rect 283389 86745 283437 86773
rect 283465 86745 283499 86773
rect 283527 86745 283561 86773
rect 283589 86745 283623 86773
rect 283651 86745 283699 86773
rect 283389 77959 283699 86745
rect 283389 77931 283437 77959
rect 283465 77931 283499 77959
rect 283527 77931 283561 77959
rect 283589 77931 283623 77959
rect 283651 77931 283699 77959
rect 283389 77897 283699 77931
rect 283389 77869 283437 77897
rect 283465 77869 283499 77897
rect 283527 77869 283561 77897
rect 283589 77869 283623 77897
rect 283651 77869 283699 77897
rect 283389 77835 283699 77869
rect 283389 77807 283437 77835
rect 283465 77807 283499 77835
rect 283527 77807 283561 77835
rect 283589 77807 283623 77835
rect 283651 77807 283699 77835
rect 283389 77773 283699 77807
rect 283389 77745 283437 77773
rect 283465 77745 283499 77773
rect 283527 77745 283561 77773
rect 283589 77745 283623 77773
rect 283651 77745 283699 77773
rect 283389 68959 283699 77745
rect 283389 68931 283437 68959
rect 283465 68931 283499 68959
rect 283527 68931 283561 68959
rect 283589 68931 283623 68959
rect 283651 68931 283699 68959
rect 283389 68897 283699 68931
rect 283389 68869 283437 68897
rect 283465 68869 283499 68897
rect 283527 68869 283561 68897
rect 283589 68869 283623 68897
rect 283651 68869 283699 68897
rect 283389 68835 283699 68869
rect 283389 68807 283437 68835
rect 283465 68807 283499 68835
rect 283527 68807 283561 68835
rect 283589 68807 283623 68835
rect 283651 68807 283699 68835
rect 283389 68773 283699 68807
rect 283389 68745 283437 68773
rect 283465 68745 283499 68773
rect 283527 68745 283561 68773
rect 283589 68745 283623 68773
rect 283651 68745 283699 68773
rect 283389 59959 283699 68745
rect 283389 59931 283437 59959
rect 283465 59931 283499 59959
rect 283527 59931 283561 59959
rect 283589 59931 283623 59959
rect 283651 59931 283699 59959
rect 283389 59897 283699 59931
rect 283389 59869 283437 59897
rect 283465 59869 283499 59897
rect 283527 59869 283561 59897
rect 283589 59869 283623 59897
rect 283651 59869 283699 59897
rect 283389 59835 283699 59869
rect 283389 59807 283437 59835
rect 283465 59807 283499 59835
rect 283527 59807 283561 59835
rect 283589 59807 283623 59835
rect 283651 59807 283699 59835
rect 283389 59773 283699 59807
rect 283389 59745 283437 59773
rect 283465 59745 283499 59773
rect 283527 59745 283561 59773
rect 283589 59745 283623 59773
rect 283651 59745 283699 59773
rect 283389 50959 283699 59745
rect 283389 50931 283437 50959
rect 283465 50931 283499 50959
rect 283527 50931 283561 50959
rect 283589 50931 283623 50959
rect 283651 50931 283699 50959
rect 283389 50897 283699 50931
rect 283389 50869 283437 50897
rect 283465 50869 283499 50897
rect 283527 50869 283561 50897
rect 283589 50869 283623 50897
rect 283651 50869 283699 50897
rect 283389 50835 283699 50869
rect 283389 50807 283437 50835
rect 283465 50807 283499 50835
rect 283527 50807 283561 50835
rect 283589 50807 283623 50835
rect 283651 50807 283699 50835
rect 283389 50773 283699 50807
rect 283389 50745 283437 50773
rect 283465 50745 283499 50773
rect 283527 50745 283561 50773
rect 283589 50745 283623 50773
rect 283651 50745 283699 50773
rect 283389 41959 283699 50745
rect 283389 41931 283437 41959
rect 283465 41931 283499 41959
rect 283527 41931 283561 41959
rect 283589 41931 283623 41959
rect 283651 41931 283699 41959
rect 283389 41897 283699 41931
rect 283389 41869 283437 41897
rect 283465 41869 283499 41897
rect 283527 41869 283561 41897
rect 283589 41869 283623 41897
rect 283651 41869 283699 41897
rect 283389 41835 283699 41869
rect 283389 41807 283437 41835
rect 283465 41807 283499 41835
rect 283527 41807 283561 41835
rect 283589 41807 283623 41835
rect 283651 41807 283699 41835
rect 283389 41773 283699 41807
rect 283389 41745 283437 41773
rect 283465 41745 283499 41773
rect 283527 41745 283561 41773
rect 283589 41745 283623 41773
rect 283651 41745 283699 41773
rect 283389 32959 283699 41745
rect 283389 32931 283437 32959
rect 283465 32931 283499 32959
rect 283527 32931 283561 32959
rect 283589 32931 283623 32959
rect 283651 32931 283699 32959
rect 283389 32897 283699 32931
rect 283389 32869 283437 32897
rect 283465 32869 283499 32897
rect 283527 32869 283561 32897
rect 283589 32869 283623 32897
rect 283651 32869 283699 32897
rect 283389 32835 283699 32869
rect 283389 32807 283437 32835
rect 283465 32807 283499 32835
rect 283527 32807 283561 32835
rect 283589 32807 283623 32835
rect 283651 32807 283699 32835
rect 283389 32773 283699 32807
rect 283389 32745 283437 32773
rect 283465 32745 283499 32773
rect 283527 32745 283561 32773
rect 283589 32745 283623 32773
rect 283651 32745 283699 32773
rect 283389 23959 283699 32745
rect 283389 23931 283437 23959
rect 283465 23931 283499 23959
rect 283527 23931 283561 23959
rect 283589 23931 283623 23959
rect 283651 23931 283699 23959
rect 283389 23897 283699 23931
rect 283389 23869 283437 23897
rect 283465 23869 283499 23897
rect 283527 23869 283561 23897
rect 283589 23869 283623 23897
rect 283651 23869 283699 23897
rect 283389 23835 283699 23869
rect 283389 23807 283437 23835
rect 283465 23807 283499 23835
rect 283527 23807 283561 23835
rect 283589 23807 283623 23835
rect 283651 23807 283699 23835
rect 283389 23773 283699 23807
rect 283389 23745 283437 23773
rect 283465 23745 283499 23773
rect 283527 23745 283561 23773
rect 283589 23745 283623 23773
rect 283651 23745 283699 23773
rect 283389 14959 283699 23745
rect 283389 14931 283437 14959
rect 283465 14931 283499 14959
rect 283527 14931 283561 14959
rect 283589 14931 283623 14959
rect 283651 14931 283699 14959
rect 283389 14897 283699 14931
rect 283389 14869 283437 14897
rect 283465 14869 283499 14897
rect 283527 14869 283561 14897
rect 283589 14869 283623 14897
rect 283651 14869 283699 14897
rect 283389 14835 283699 14869
rect 283389 14807 283437 14835
rect 283465 14807 283499 14835
rect 283527 14807 283561 14835
rect 283589 14807 283623 14835
rect 283651 14807 283699 14835
rect 283389 14773 283699 14807
rect 283389 14745 283437 14773
rect 283465 14745 283499 14773
rect 283527 14745 283561 14773
rect 283589 14745 283623 14773
rect 283651 14745 283699 14773
rect 283389 5959 283699 14745
rect 283389 5931 283437 5959
rect 283465 5931 283499 5959
rect 283527 5931 283561 5959
rect 283589 5931 283623 5959
rect 283651 5931 283699 5959
rect 283389 5897 283699 5931
rect 283389 5869 283437 5897
rect 283465 5869 283499 5897
rect 283527 5869 283561 5897
rect 283589 5869 283623 5897
rect 283651 5869 283699 5897
rect 283389 5835 283699 5869
rect 283389 5807 283437 5835
rect 283465 5807 283499 5835
rect 283527 5807 283561 5835
rect 283589 5807 283623 5835
rect 283651 5807 283699 5835
rect 283389 5773 283699 5807
rect 283389 5745 283437 5773
rect 283465 5745 283499 5773
rect 283527 5745 283561 5773
rect 283589 5745 283623 5773
rect 283651 5745 283699 5773
rect 283389 424 283699 5745
rect 283389 396 283437 424
rect 283465 396 283499 424
rect 283527 396 283561 424
rect 283589 396 283623 424
rect 283651 396 283699 424
rect 283389 362 283699 396
rect 283389 334 283437 362
rect 283465 334 283499 362
rect 283527 334 283561 362
rect 283589 334 283623 362
rect 283651 334 283699 362
rect 283389 300 283699 334
rect 283389 272 283437 300
rect 283465 272 283499 300
rect 283527 272 283561 300
rect 283589 272 283623 300
rect 283651 272 283699 300
rect 283389 238 283699 272
rect 283389 210 283437 238
rect 283465 210 283499 238
rect 283527 210 283561 238
rect 283589 210 283623 238
rect 283651 210 283699 238
rect 283389 162 283699 210
rect 290529 299190 290839 299718
rect 290529 299162 290577 299190
rect 290605 299162 290639 299190
rect 290667 299162 290701 299190
rect 290729 299162 290763 299190
rect 290791 299162 290839 299190
rect 290529 299128 290839 299162
rect 290529 299100 290577 299128
rect 290605 299100 290639 299128
rect 290667 299100 290701 299128
rect 290729 299100 290763 299128
rect 290791 299100 290839 299128
rect 290529 299066 290839 299100
rect 290529 299038 290577 299066
rect 290605 299038 290639 299066
rect 290667 299038 290701 299066
rect 290729 299038 290763 299066
rect 290791 299038 290839 299066
rect 290529 299004 290839 299038
rect 290529 298976 290577 299004
rect 290605 298976 290639 299004
rect 290667 298976 290701 299004
rect 290729 298976 290763 299004
rect 290791 298976 290839 299004
rect 290529 290959 290839 298976
rect 290529 290931 290577 290959
rect 290605 290931 290639 290959
rect 290667 290931 290701 290959
rect 290729 290931 290763 290959
rect 290791 290931 290839 290959
rect 290529 290897 290839 290931
rect 290529 290869 290577 290897
rect 290605 290869 290639 290897
rect 290667 290869 290701 290897
rect 290729 290869 290763 290897
rect 290791 290869 290839 290897
rect 290529 290835 290839 290869
rect 290529 290807 290577 290835
rect 290605 290807 290639 290835
rect 290667 290807 290701 290835
rect 290729 290807 290763 290835
rect 290791 290807 290839 290835
rect 290529 290773 290839 290807
rect 290529 290745 290577 290773
rect 290605 290745 290639 290773
rect 290667 290745 290701 290773
rect 290729 290745 290763 290773
rect 290791 290745 290839 290773
rect 290529 281959 290839 290745
rect 290529 281931 290577 281959
rect 290605 281931 290639 281959
rect 290667 281931 290701 281959
rect 290729 281931 290763 281959
rect 290791 281931 290839 281959
rect 290529 281897 290839 281931
rect 290529 281869 290577 281897
rect 290605 281869 290639 281897
rect 290667 281869 290701 281897
rect 290729 281869 290763 281897
rect 290791 281869 290839 281897
rect 290529 281835 290839 281869
rect 290529 281807 290577 281835
rect 290605 281807 290639 281835
rect 290667 281807 290701 281835
rect 290729 281807 290763 281835
rect 290791 281807 290839 281835
rect 290529 281773 290839 281807
rect 290529 281745 290577 281773
rect 290605 281745 290639 281773
rect 290667 281745 290701 281773
rect 290729 281745 290763 281773
rect 290791 281745 290839 281773
rect 290529 272959 290839 281745
rect 290529 272931 290577 272959
rect 290605 272931 290639 272959
rect 290667 272931 290701 272959
rect 290729 272931 290763 272959
rect 290791 272931 290839 272959
rect 290529 272897 290839 272931
rect 290529 272869 290577 272897
rect 290605 272869 290639 272897
rect 290667 272869 290701 272897
rect 290729 272869 290763 272897
rect 290791 272869 290839 272897
rect 290529 272835 290839 272869
rect 290529 272807 290577 272835
rect 290605 272807 290639 272835
rect 290667 272807 290701 272835
rect 290729 272807 290763 272835
rect 290791 272807 290839 272835
rect 290529 272773 290839 272807
rect 290529 272745 290577 272773
rect 290605 272745 290639 272773
rect 290667 272745 290701 272773
rect 290729 272745 290763 272773
rect 290791 272745 290839 272773
rect 290529 263959 290839 272745
rect 290529 263931 290577 263959
rect 290605 263931 290639 263959
rect 290667 263931 290701 263959
rect 290729 263931 290763 263959
rect 290791 263931 290839 263959
rect 290529 263897 290839 263931
rect 290529 263869 290577 263897
rect 290605 263869 290639 263897
rect 290667 263869 290701 263897
rect 290729 263869 290763 263897
rect 290791 263869 290839 263897
rect 290529 263835 290839 263869
rect 290529 263807 290577 263835
rect 290605 263807 290639 263835
rect 290667 263807 290701 263835
rect 290729 263807 290763 263835
rect 290791 263807 290839 263835
rect 290529 263773 290839 263807
rect 290529 263745 290577 263773
rect 290605 263745 290639 263773
rect 290667 263745 290701 263773
rect 290729 263745 290763 263773
rect 290791 263745 290839 263773
rect 290529 254959 290839 263745
rect 290529 254931 290577 254959
rect 290605 254931 290639 254959
rect 290667 254931 290701 254959
rect 290729 254931 290763 254959
rect 290791 254931 290839 254959
rect 290529 254897 290839 254931
rect 290529 254869 290577 254897
rect 290605 254869 290639 254897
rect 290667 254869 290701 254897
rect 290729 254869 290763 254897
rect 290791 254869 290839 254897
rect 290529 254835 290839 254869
rect 290529 254807 290577 254835
rect 290605 254807 290639 254835
rect 290667 254807 290701 254835
rect 290729 254807 290763 254835
rect 290791 254807 290839 254835
rect 290529 254773 290839 254807
rect 290529 254745 290577 254773
rect 290605 254745 290639 254773
rect 290667 254745 290701 254773
rect 290729 254745 290763 254773
rect 290791 254745 290839 254773
rect 290529 245959 290839 254745
rect 290529 245931 290577 245959
rect 290605 245931 290639 245959
rect 290667 245931 290701 245959
rect 290729 245931 290763 245959
rect 290791 245931 290839 245959
rect 290529 245897 290839 245931
rect 290529 245869 290577 245897
rect 290605 245869 290639 245897
rect 290667 245869 290701 245897
rect 290729 245869 290763 245897
rect 290791 245869 290839 245897
rect 290529 245835 290839 245869
rect 290529 245807 290577 245835
rect 290605 245807 290639 245835
rect 290667 245807 290701 245835
rect 290729 245807 290763 245835
rect 290791 245807 290839 245835
rect 290529 245773 290839 245807
rect 290529 245745 290577 245773
rect 290605 245745 290639 245773
rect 290667 245745 290701 245773
rect 290729 245745 290763 245773
rect 290791 245745 290839 245773
rect 290529 236959 290839 245745
rect 290529 236931 290577 236959
rect 290605 236931 290639 236959
rect 290667 236931 290701 236959
rect 290729 236931 290763 236959
rect 290791 236931 290839 236959
rect 290529 236897 290839 236931
rect 290529 236869 290577 236897
rect 290605 236869 290639 236897
rect 290667 236869 290701 236897
rect 290729 236869 290763 236897
rect 290791 236869 290839 236897
rect 290529 236835 290839 236869
rect 290529 236807 290577 236835
rect 290605 236807 290639 236835
rect 290667 236807 290701 236835
rect 290729 236807 290763 236835
rect 290791 236807 290839 236835
rect 290529 236773 290839 236807
rect 290529 236745 290577 236773
rect 290605 236745 290639 236773
rect 290667 236745 290701 236773
rect 290729 236745 290763 236773
rect 290791 236745 290839 236773
rect 290529 227959 290839 236745
rect 290529 227931 290577 227959
rect 290605 227931 290639 227959
rect 290667 227931 290701 227959
rect 290729 227931 290763 227959
rect 290791 227931 290839 227959
rect 290529 227897 290839 227931
rect 290529 227869 290577 227897
rect 290605 227869 290639 227897
rect 290667 227869 290701 227897
rect 290729 227869 290763 227897
rect 290791 227869 290839 227897
rect 290529 227835 290839 227869
rect 290529 227807 290577 227835
rect 290605 227807 290639 227835
rect 290667 227807 290701 227835
rect 290729 227807 290763 227835
rect 290791 227807 290839 227835
rect 290529 227773 290839 227807
rect 290529 227745 290577 227773
rect 290605 227745 290639 227773
rect 290667 227745 290701 227773
rect 290729 227745 290763 227773
rect 290791 227745 290839 227773
rect 290529 218959 290839 227745
rect 290529 218931 290577 218959
rect 290605 218931 290639 218959
rect 290667 218931 290701 218959
rect 290729 218931 290763 218959
rect 290791 218931 290839 218959
rect 290529 218897 290839 218931
rect 290529 218869 290577 218897
rect 290605 218869 290639 218897
rect 290667 218869 290701 218897
rect 290729 218869 290763 218897
rect 290791 218869 290839 218897
rect 290529 218835 290839 218869
rect 290529 218807 290577 218835
rect 290605 218807 290639 218835
rect 290667 218807 290701 218835
rect 290729 218807 290763 218835
rect 290791 218807 290839 218835
rect 290529 218773 290839 218807
rect 290529 218745 290577 218773
rect 290605 218745 290639 218773
rect 290667 218745 290701 218773
rect 290729 218745 290763 218773
rect 290791 218745 290839 218773
rect 290529 209959 290839 218745
rect 290529 209931 290577 209959
rect 290605 209931 290639 209959
rect 290667 209931 290701 209959
rect 290729 209931 290763 209959
rect 290791 209931 290839 209959
rect 290529 209897 290839 209931
rect 290529 209869 290577 209897
rect 290605 209869 290639 209897
rect 290667 209869 290701 209897
rect 290729 209869 290763 209897
rect 290791 209869 290839 209897
rect 290529 209835 290839 209869
rect 290529 209807 290577 209835
rect 290605 209807 290639 209835
rect 290667 209807 290701 209835
rect 290729 209807 290763 209835
rect 290791 209807 290839 209835
rect 290529 209773 290839 209807
rect 290529 209745 290577 209773
rect 290605 209745 290639 209773
rect 290667 209745 290701 209773
rect 290729 209745 290763 209773
rect 290791 209745 290839 209773
rect 290529 200959 290839 209745
rect 290529 200931 290577 200959
rect 290605 200931 290639 200959
rect 290667 200931 290701 200959
rect 290729 200931 290763 200959
rect 290791 200931 290839 200959
rect 290529 200897 290839 200931
rect 290529 200869 290577 200897
rect 290605 200869 290639 200897
rect 290667 200869 290701 200897
rect 290729 200869 290763 200897
rect 290791 200869 290839 200897
rect 290529 200835 290839 200869
rect 290529 200807 290577 200835
rect 290605 200807 290639 200835
rect 290667 200807 290701 200835
rect 290729 200807 290763 200835
rect 290791 200807 290839 200835
rect 290529 200773 290839 200807
rect 290529 200745 290577 200773
rect 290605 200745 290639 200773
rect 290667 200745 290701 200773
rect 290729 200745 290763 200773
rect 290791 200745 290839 200773
rect 290529 191959 290839 200745
rect 290529 191931 290577 191959
rect 290605 191931 290639 191959
rect 290667 191931 290701 191959
rect 290729 191931 290763 191959
rect 290791 191931 290839 191959
rect 290529 191897 290839 191931
rect 290529 191869 290577 191897
rect 290605 191869 290639 191897
rect 290667 191869 290701 191897
rect 290729 191869 290763 191897
rect 290791 191869 290839 191897
rect 290529 191835 290839 191869
rect 290529 191807 290577 191835
rect 290605 191807 290639 191835
rect 290667 191807 290701 191835
rect 290729 191807 290763 191835
rect 290791 191807 290839 191835
rect 290529 191773 290839 191807
rect 290529 191745 290577 191773
rect 290605 191745 290639 191773
rect 290667 191745 290701 191773
rect 290729 191745 290763 191773
rect 290791 191745 290839 191773
rect 290529 182959 290839 191745
rect 290529 182931 290577 182959
rect 290605 182931 290639 182959
rect 290667 182931 290701 182959
rect 290729 182931 290763 182959
rect 290791 182931 290839 182959
rect 290529 182897 290839 182931
rect 290529 182869 290577 182897
rect 290605 182869 290639 182897
rect 290667 182869 290701 182897
rect 290729 182869 290763 182897
rect 290791 182869 290839 182897
rect 290529 182835 290839 182869
rect 290529 182807 290577 182835
rect 290605 182807 290639 182835
rect 290667 182807 290701 182835
rect 290729 182807 290763 182835
rect 290791 182807 290839 182835
rect 290529 182773 290839 182807
rect 290529 182745 290577 182773
rect 290605 182745 290639 182773
rect 290667 182745 290701 182773
rect 290729 182745 290763 182773
rect 290791 182745 290839 182773
rect 290529 173959 290839 182745
rect 290529 173931 290577 173959
rect 290605 173931 290639 173959
rect 290667 173931 290701 173959
rect 290729 173931 290763 173959
rect 290791 173931 290839 173959
rect 290529 173897 290839 173931
rect 290529 173869 290577 173897
rect 290605 173869 290639 173897
rect 290667 173869 290701 173897
rect 290729 173869 290763 173897
rect 290791 173869 290839 173897
rect 290529 173835 290839 173869
rect 290529 173807 290577 173835
rect 290605 173807 290639 173835
rect 290667 173807 290701 173835
rect 290729 173807 290763 173835
rect 290791 173807 290839 173835
rect 290529 173773 290839 173807
rect 290529 173745 290577 173773
rect 290605 173745 290639 173773
rect 290667 173745 290701 173773
rect 290729 173745 290763 173773
rect 290791 173745 290839 173773
rect 290529 164959 290839 173745
rect 290529 164931 290577 164959
rect 290605 164931 290639 164959
rect 290667 164931 290701 164959
rect 290729 164931 290763 164959
rect 290791 164931 290839 164959
rect 290529 164897 290839 164931
rect 290529 164869 290577 164897
rect 290605 164869 290639 164897
rect 290667 164869 290701 164897
rect 290729 164869 290763 164897
rect 290791 164869 290839 164897
rect 290529 164835 290839 164869
rect 290529 164807 290577 164835
rect 290605 164807 290639 164835
rect 290667 164807 290701 164835
rect 290729 164807 290763 164835
rect 290791 164807 290839 164835
rect 290529 164773 290839 164807
rect 290529 164745 290577 164773
rect 290605 164745 290639 164773
rect 290667 164745 290701 164773
rect 290729 164745 290763 164773
rect 290791 164745 290839 164773
rect 290529 155959 290839 164745
rect 290529 155931 290577 155959
rect 290605 155931 290639 155959
rect 290667 155931 290701 155959
rect 290729 155931 290763 155959
rect 290791 155931 290839 155959
rect 290529 155897 290839 155931
rect 290529 155869 290577 155897
rect 290605 155869 290639 155897
rect 290667 155869 290701 155897
rect 290729 155869 290763 155897
rect 290791 155869 290839 155897
rect 290529 155835 290839 155869
rect 290529 155807 290577 155835
rect 290605 155807 290639 155835
rect 290667 155807 290701 155835
rect 290729 155807 290763 155835
rect 290791 155807 290839 155835
rect 290529 155773 290839 155807
rect 290529 155745 290577 155773
rect 290605 155745 290639 155773
rect 290667 155745 290701 155773
rect 290729 155745 290763 155773
rect 290791 155745 290839 155773
rect 290529 146959 290839 155745
rect 290529 146931 290577 146959
rect 290605 146931 290639 146959
rect 290667 146931 290701 146959
rect 290729 146931 290763 146959
rect 290791 146931 290839 146959
rect 290529 146897 290839 146931
rect 290529 146869 290577 146897
rect 290605 146869 290639 146897
rect 290667 146869 290701 146897
rect 290729 146869 290763 146897
rect 290791 146869 290839 146897
rect 290529 146835 290839 146869
rect 290529 146807 290577 146835
rect 290605 146807 290639 146835
rect 290667 146807 290701 146835
rect 290729 146807 290763 146835
rect 290791 146807 290839 146835
rect 290529 146773 290839 146807
rect 290529 146745 290577 146773
rect 290605 146745 290639 146773
rect 290667 146745 290701 146773
rect 290729 146745 290763 146773
rect 290791 146745 290839 146773
rect 290529 137959 290839 146745
rect 290529 137931 290577 137959
rect 290605 137931 290639 137959
rect 290667 137931 290701 137959
rect 290729 137931 290763 137959
rect 290791 137931 290839 137959
rect 290529 137897 290839 137931
rect 290529 137869 290577 137897
rect 290605 137869 290639 137897
rect 290667 137869 290701 137897
rect 290729 137869 290763 137897
rect 290791 137869 290839 137897
rect 290529 137835 290839 137869
rect 290529 137807 290577 137835
rect 290605 137807 290639 137835
rect 290667 137807 290701 137835
rect 290729 137807 290763 137835
rect 290791 137807 290839 137835
rect 290529 137773 290839 137807
rect 290529 137745 290577 137773
rect 290605 137745 290639 137773
rect 290667 137745 290701 137773
rect 290729 137745 290763 137773
rect 290791 137745 290839 137773
rect 290529 128959 290839 137745
rect 290529 128931 290577 128959
rect 290605 128931 290639 128959
rect 290667 128931 290701 128959
rect 290729 128931 290763 128959
rect 290791 128931 290839 128959
rect 290529 128897 290839 128931
rect 290529 128869 290577 128897
rect 290605 128869 290639 128897
rect 290667 128869 290701 128897
rect 290729 128869 290763 128897
rect 290791 128869 290839 128897
rect 290529 128835 290839 128869
rect 290529 128807 290577 128835
rect 290605 128807 290639 128835
rect 290667 128807 290701 128835
rect 290729 128807 290763 128835
rect 290791 128807 290839 128835
rect 290529 128773 290839 128807
rect 290529 128745 290577 128773
rect 290605 128745 290639 128773
rect 290667 128745 290701 128773
rect 290729 128745 290763 128773
rect 290791 128745 290839 128773
rect 290529 119959 290839 128745
rect 290529 119931 290577 119959
rect 290605 119931 290639 119959
rect 290667 119931 290701 119959
rect 290729 119931 290763 119959
rect 290791 119931 290839 119959
rect 290529 119897 290839 119931
rect 290529 119869 290577 119897
rect 290605 119869 290639 119897
rect 290667 119869 290701 119897
rect 290729 119869 290763 119897
rect 290791 119869 290839 119897
rect 290529 119835 290839 119869
rect 290529 119807 290577 119835
rect 290605 119807 290639 119835
rect 290667 119807 290701 119835
rect 290729 119807 290763 119835
rect 290791 119807 290839 119835
rect 290529 119773 290839 119807
rect 290529 119745 290577 119773
rect 290605 119745 290639 119773
rect 290667 119745 290701 119773
rect 290729 119745 290763 119773
rect 290791 119745 290839 119773
rect 290529 110959 290839 119745
rect 290529 110931 290577 110959
rect 290605 110931 290639 110959
rect 290667 110931 290701 110959
rect 290729 110931 290763 110959
rect 290791 110931 290839 110959
rect 290529 110897 290839 110931
rect 290529 110869 290577 110897
rect 290605 110869 290639 110897
rect 290667 110869 290701 110897
rect 290729 110869 290763 110897
rect 290791 110869 290839 110897
rect 290529 110835 290839 110869
rect 290529 110807 290577 110835
rect 290605 110807 290639 110835
rect 290667 110807 290701 110835
rect 290729 110807 290763 110835
rect 290791 110807 290839 110835
rect 290529 110773 290839 110807
rect 290529 110745 290577 110773
rect 290605 110745 290639 110773
rect 290667 110745 290701 110773
rect 290729 110745 290763 110773
rect 290791 110745 290839 110773
rect 290529 101959 290839 110745
rect 290529 101931 290577 101959
rect 290605 101931 290639 101959
rect 290667 101931 290701 101959
rect 290729 101931 290763 101959
rect 290791 101931 290839 101959
rect 290529 101897 290839 101931
rect 290529 101869 290577 101897
rect 290605 101869 290639 101897
rect 290667 101869 290701 101897
rect 290729 101869 290763 101897
rect 290791 101869 290839 101897
rect 290529 101835 290839 101869
rect 290529 101807 290577 101835
rect 290605 101807 290639 101835
rect 290667 101807 290701 101835
rect 290729 101807 290763 101835
rect 290791 101807 290839 101835
rect 290529 101773 290839 101807
rect 290529 101745 290577 101773
rect 290605 101745 290639 101773
rect 290667 101745 290701 101773
rect 290729 101745 290763 101773
rect 290791 101745 290839 101773
rect 290529 92959 290839 101745
rect 290529 92931 290577 92959
rect 290605 92931 290639 92959
rect 290667 92931 290701 92959
rect 290729 92931 290763 92959
rect 290791 92931 290839 92959
rect 290529 92897 290839 92931
rect 290529 92869 290577 92897
rect 290605 92869 290639 92897
rect 290667 92869 290701 92897
rect 290729 92869 290763 92897
rect 290791 92869 290839 92897
rect 290529 92835 290839 92869
rect 290529 92807 290577 92835
rect 290605 92807 290639 92835
rect 290667 92807 290701 92835
rect 290729 92807 290763 92835
rect 290791 92807 290839 92835
rect 290529 92773 290839 92807
rect 290529 92745 290577 92773
rect 290605 92745 290639 92773
rect 290667 92745 290701 92773
rect 290729 92745 290763 92773
rect 290791 92745 290839 92773
rect 290529 83959 290839 92745
rect 290529 83931 290577 83959
rect 290605 83931 290639 83959
rect 290667 83931 290701 83959
rect 290729 83931 290763 83959
rect 290791 83931 290839 83959
rect 290529 83897 290839 83931
rect 290529 83869 290577 83897
rect 290605 83869 290639 83897
rect 290667 83869 290701 83897
rect 290729 83869 290763 83897
rect 290791 83869 290839 83897
rect 290529 83835 290839 83869
rect 290529 83807 290577 83835
rect 290605 83807 290639 83835
rect 290667 83807 290701 83835
rect 290729 83807 290763 83835
rect 290791 83807 290839 83835
rect 290529 83773 290839 83807
rect 290529 83745 290577 83773
rect 290605 83745 290639 83773
rect 290667 83745 290701 83773
rect 290729 83745 290763 83773
rect 290791 83745 290839 83773
rect 290529 74959 290839 83745
rect 290529 74931 290577 74959
rect 290605 74931 290639 74959
rect 290667 74931 290701 74959
rect 290729 74931 290763 74959
rect 290791 74931 290839 74959
rect 290529 74897 290839 74931
rect 290529 74869 290577 74897
rect 290605 74869 290639 74897
rect 290667 74869 290701 74897
rect 290729 74869 290763 74897
rect 290791 74869 290839 74897
rect 290529 74835 290839 74869
rect 290529 74807 290577 74835
rect 290605 74807 290639 74835
rect 290667 74807 290701 74835
rect 290729 74807 290763 74835
rect 290791 74807 290839 74835
rect 290529 74773 290839 74807
rect 290529 74745 290577 74773
rect 290605 74745 290639 74773
rect 290667 74745 290701 74773
rect 290729 74745 290763 74773
rect 290791 74745 290839 74773
rect 290529 65959 290839 74745
rect 290529 65931 290577 65959
rect 290605 65931 290639 65959
rect 290667 65931 290701 65959
rect 290729 65931 290763 65959
rect 290791 65931 290839 65959
rect 290529 65897 290839 65931
rect 290529 65869 290577 65897
rect 290605 65869 290639 65897
rect 290667 65869 290701 65897
rect 290729 65869 290763 65897
rect 290791 65869 290839 65897
rect 290529 65835 290839 65869
rect 290529 65807 290577 65835
rect 290605 65807 290639 65835
rect 290667 65807 290701 65835
rect 290729 65807 290763 65835
rect 290791 65807 290839 65835
rect 290529 65773 290839 65807
rect 290529 65745 290577 65773
rect 290605 65745 290639 65773
rect 290667 65745 290701 65773
rect 290729 65745 290763 65773
rect 290791 65745 290839 65773
rect 290529 56959 290839 65745
rect 290529 56931 290577 56959
rect 290605 56931 290639 56959
rect 290667 56931 290701 56959
rect 290729 56931 290763 56959
rect 290791 56931 290839 56959
rect 290529 56897 290839 56931
rect 290529 56869 290577 56897
rect 290605 56869 290639 56897
rect 290667 56869 290701 56897
rect 290729 56869 290763 56897
rect 290791 56869 290839 56897
rect 290529 56835 290839 56869
rect 290529 56807 290577 56835
rect 290605 56807 290639 56835
rect 290667 56807 290701 56835
rect 290729 56807 290763 56835
rect 290791 56807 290839 56835
rect 290529 56773 290839 56807
rect 290529 56745 290577 56773
rect 290605 56745 290639 56773
rect 290667 56745 290701 56773
rect 290729 56745 290763 56773
rect 290791 56745 290839 56773
rect 290529 47959 290839 56745
rect 290529 47931 290577 47959
rect 290605 47931 290639 47959
rect 290667 47931 290701 47959
rect 290729 47931 290763 47959
rect 290791 47931 290839 47959
rect 290529 47897 290839 47931
rect 290529 47869 290577 47897
rect 290605 47869 290639 47897
rect 290667 47869 290701 47897
rect 290729 47869 290763 47897
rect 290791 47869 290839 47897
rect 290529 47835 290839 47869
rect 290529 47807 290577 47835
rect 290605 47807 290639 47835
rect 290667 47807 290701 47835
rect 290729 47807 290763 47835
rect 290791 47807 290839 47835
rect 290529 47773 290839 47807
rect 290529 47745 290577 47773
rect 290605 47745 290639 47773
rect 290667 47745 290701 47773
rect 290729 47745 290763 47773
rect 290791 47745 290839 47773
rect 290529 38959 290839 47745
rect 290529 38931 290577 38959
rect 290605 38931 290639 38959
rect 290667 38931 290701 38959
rect 290729 38931 290763 38959
rect 290791 38931 290839 38959
rect 290529 38897 290839 38931
rect 290529 38869 290577 38897
rect 290605 38869 290639 38897
rect 290667 38869 290701 38897
rect 290729 38869 290763 38897
rect 290791 38869 290839 38897
rect 290529 38835 290839 38869
rect 290529 38807 290577 38835
rect 290605 38807 290639 38835
rect 290667 38807 290701 38835
rect 290729 38807 290763 38835
rect 290791 38807 290839 38835
rect 290529 38773 290839 38807
rect 290529 38745 290577 38773
rect 290605 38745 290639 38773
rect 290667 38745 290701 38773
rect 290729 38745 290763 38773
rect 290791 38745 290839 38773
rect 290529 29959 290839 38745
rect 290529 29931 290577 29959
rect 290605 29931 290639 29959
rect 290667 29931 290701 29959
rect 290729 29931 290763 29959
rect 290791 29931 290839 29959
rect 290529 29897 290839 29931
rect 290529 29869 290577 29897
rect 290605 29869 290639 29897
rect 290667 29869 290701 29897
rect 290729 29869 290763 29897
rect 290791 29869 290839 29897
rect 290529 29835 290839 29869
rect 290529 29807 290577 29835
rect 290605 29807 290639 29835
rect 290667 29807 290701 29835
rect 290729 29807 290763 29835
rect 290791 29807 290839 29835
rect 290529 29773 290839 29807
rect 290529 29745 290577 29773
rect 290605 29745 290639 29773
rect 290667 29745 290701 29773
rect 290729 29745 290763 29773
rect 290791 29745 290839 29773
rect 290529 20959 290839 29745
rect 290529 20931 290577 20959
rect 290605 20931 290639 20959
rect 290667 20931 290701 20959
rect 290729 20931 290763 20959
rect 290791 20931 290839 20959
rect 290529 20897 290839 20931
rect 290529 20869 290577 20897
rect 290605 20869 290639 20897
rect 290667 20869 290701 20897
rect 290729 20869 290763 20897
rect 290791 20869 290839 20897
rect 290529 20835 290839 20869
rect 290529 20807 290577 20835
rect 290605 20807 290639 20835
rect 290667 20807 290701 20835
rect 290729 20807 290763 20835
rect 290791 20807 290839 20835
rect 290529 20773 290839 20807
rect 290529 20745 290577 20773
rect 290605 20745 290639 20773
rect 290667 20745 290701 20773
rect 290729 20745 290763 20773
rect 290791 20745 290839 20773
rect 290529 11959 290839 20745
rect 290529 11931 290577 11959
rect 290605 11931 290639 11959
rect 290667 11931 290701 11959
rect 290729 11931 290763 11959
rect 290791 11931 290839 11959
rect 290529 11897 290839 11931
rect 290529 11869 290577 11897
rect 290605 11869 290639 11897
rect 290667 11869 290701 11897
rect 290729 11869 290763 11897
rect 290791 11869 290839 11897
rect 290529 11835 290839 11869
rect 290529 11807 290577 11835
rect 290605 11807 290639 11835
rect 290667 11807 290701 11835
rect 290729 11807 290763 11835
rect 290791 11807 290839 11835
rect 290529 11773 290839 11807
rect 290529 11745 290577 11773
rect 290605 11745 290639 11773
rect 290667 11745 290701 11773
rect 290729 11745 290763 11773
rect 290791 11745 290839 11773
rect 290529 2959 290839 11745
rect 290529 2931 290577 2959
rect 290605 2931 290639 2959
rect 290667 2931 290701 2959
rect 290729 2931 290763 2959
rect 290791 2931 290839 2959
rect 290529 2897 290839 2931
rect 290529 2869 290577 2897
rect 290605 2869 290639 2897
rect 290667 2869 290701 2897
rect 290729 2869 290763 2897
rect 290791 2869 290839 2897
rect 290529 2835 290839 2869
rect 290529 2807 290577 2835
rect 290605 2807 290639 2835
rect 290667 2807 290701 2835
rect 290729 2807 290763 2835
rect 290791 2807 290839 2835
rect 290529 2773 290839 2807
rect 290529 2745 290577 2773
rect 290605 2745 290639 2773
rect 290667 2745 290701 2773
rect 290729 2745 290763 2773
rect 290791 2745 290839 2773
rect 290529 904 290839 2745
rect 290529 876 290577 904
rect 290605 876 290639 904
rect 290667 876 290701 904
rect 290729 876 290763 904
rect 290791 876 290839 904
rect 290529 842 290839 876
rect 290529 814 290577 842
rect 290605 814 290639 842
rect 290667 814 290701 842
rect 290729 814 290763 842
rect 290791 814 290839 842
rect 290529 780 290839 814
rect 290529 752 290577 780
rect 290605 752 290639 780
rect 290667 752 290701 780
rect 290729 752 290763 780
rect 290791 752 290839 780
rect 290529 718 290839 752
rect 290529 690 290577 718
rect 290605 690 290639 718
rect 290667 690 290701 718
rect 290729 690 290763 718
rect 290791 690 290839 718
rect 290529 162 290839 690
rect 292389 299670 292699 299718
rect 292389 299642 292437 299670
rect 292465 299642 292499 299670
rect 292527 299642 292561 299670
rect 292589 299642 292623 299670
rect 292651 299642 292699 299670
rect 292389 299608 292699 299642
rect 292389 299580 292437 299608
rect 292465 299580 292499 299608
rect 292527 299580 292561 299608
rect 292589 299580 292623 299608
rect 292651 299580 292699 299608
rect 292389 299546 292699 299580
rect 292389 299518 292437 299546
rect 292465 299518 292499 299546
rect 292527 299518 292561 299546
rect 292589 299518 292623 299546
rect 292651 299518 292699 299546
rect 292389 299484 292699 299518
rect 292389 299456 292437 299484
rect 292465 299456 292499 299484
rect 292527 299456 292561 299484
rect 292589 299456 292623 299484
rect 292651 299456 292699 299484
rect 292389 293959 292699 299456
rect 299688 299670 299998 299718
rect 299688 299642 299736 299670
rect 299764 299642 299798 299670
rect 299826 299642 299860 299670
rect 299888 299642 299922 299670
rect 299950 299642 299998 299670
rect 299688 299608 299998 299642
rect 299688 299580 299736 299608
rect 299764 299580 299798 299608
rect 299826 299580 299860 299608
rect 299888 299580 299922 299608
rect 299950 299580 299998 299608
rect 299688 299546 299998 299580
rect 299688 299518 299736 299546
rect 299764 299518 299798 299546
rect 299826 299518 299860 299546
rect 299888 299518 299922 299546
rect 299950 299518 299998 299546
rect 299688 299484 299998 299518
rect 299688 299456 299736 299484
rect 299764 299456 299798 299484
rect 299826 299456 299860 299484
rect 299888 299456 299922 299484
rect 299950 299456 299998 299484
rect 292389 293931 292437 293959
rect 292465 293931 292499 293959
rect 292527 293931 292561 293959
rect 292589 293931 292623 293959
rect 292651 293931 292699 293959
rect 292389 293897 292699 293931
rect 292389 293869 292437 293897
rect 292465 293869 292499 293897
rect 292527 293869 292561 293897
rect 292589 293869 292623 293897
rect 292651 293869 292699 293897
rect 292389 293835 292699 293869
rect 292389 293807 292437 293835
rect 292465 293807 292499 293835
rect 292527 293807 292561 293835
rect 292589 293807 292623 293835
rect 292651 293807 292699 293835
rect 292389 293773 292699 293807
rect 292389 293745 292437 293773
rect 292465 293745 292499 293773
rect 292527 293745 292561 293773
rect 292589 293745 292623 293773
rect 292651 293745 292699 293773
rect 292389 284959 292699 293745
rect 292389 284931 292437 284959
rect 292465 284931 292499 284959
rect 292527 284931 292561 284959
rect 292589 284931 292623 284959
rect 292651 284931 292699 284959
rect 292389 284897 292699 284931
rect 292389 284869 292437 284897
rect 292465 284869 292499 284897
rect 292527 284869 292561 284897
rect 292589 284869 292623 284897
rect 292651 284869 292699 284897
rect 292389 284835 292699 284869
rect 292389 284807 292437 284835
rect 292465 284807 292499 284835
rect 292527 284807 292561 284835
rect 292589 284807 292623 284835
rect 292651 284807 292699 284835
rect 292389 284773 292699 284807
rect 292389 284745 292437 284773
rect 292465 284745 292499 284773
rect 292527 284745 292561 284773
rect 292589 284745 292623 284773
rect 292651 284745 292699 284773
rect 292389 275959 292699 284745
rect 292389 275931 292437 275959
rect 292465 275931 292499 275959
rect 292527 275931 292561 275959
rect 292589 275931 292623 275959
rect 292651 275931 292699 275959
rect 292389 275897 292699 275931
rect 292389 275869 292437 275897
rect 292465 275869 292499 275897
rect 292527 275869 292561 275897
rect 292589 275869 292623 275897
rect 292651 275869 292699 275897
rect 292389 275835 292699 275869
rect 292389 275807 292437 275835
rect 292465 275807 292499 275835
rect 292527 275807 292561 275835
rect 292589 275807 292623 275835
rect 292651 275807 292699 275835
rect 292389 275773 292699 275807
rect 292389 275745 292437 275773
rect 292465 275745 292499 275773
rect 292527 275745 292561 275773
rect 292589 275745 292623 275773
rect 292651 275745 292699 275773
rect 292389 266959 292699 275745
rect 292389 266931 292437 266959
rect 292465 266931 292499 266959
rect 292527 266931 292561 266959
rect 292589 266931 292623 266959
rect 292651 266931 292699 266959
rect 292389 266897 292699 266931
rect 292389 266869 292437 266897
rect 292465 266869 292499 266897
rect 292527 266869 292561 266897
rect 292589 266869 292623 266897
rect 292651 266869 292699 266897
rect 292389 266835 292699 266869
rect 292389 266807 292437 266835
rect 292465 266807 292499 266835
rect 292527 266807 292561 266835
rect 292589 266807 292623 266835
rect 292651 266807 292699 266835
rect 292389 266773 292699 266807
rect 292389 266745 292437 266773
rect 292465 266745 292499 266773
rect 292527 266745 292561 266773
rect 292589 266745 292623 266773
rect 292651 266745 292699 266773
rect 292389 257959 292699 266745
rect 292389 257931 292437 257959
rect 292465 257931 292499 257959
rect 292527 257931 292561 257959
rect 292589 257931 292623 257959
rect 292651 257931 292699 257959
rect 292389 257897 292699 257931
rect 292389 257869 292437 257897
rect 292465 257869 292499 257897
rect 292527 257869 292561 257897
rect 292589 257869 292623 257897
rect 292651 257869 292699 257897
rect 292389 257835 292699 257869
rect 292389 257807 292437 257835
rect 292465 257807 292499 257835
rect 292527 257807 292561 257835
rect 292589 257807 292623 257835
rect 292651 257807 292699 257835
rect 292389 257773 292699 257807
rect 292389 257745 292437 257773
rect 292465 257745 292499 257773
rect 292527 257745 292561 257773
rect 292589 257745 292623 257773
rect 292651 257745 292699 257773
rect 292389 248959 292699 257745
rect 292389 248931 292437 248959
rect 292465 248931 292499 248959
rect 292527 248931 292561 248959
rect 292589 248931 292623 248959
rect 292651 248931 292699 248959
rect 292389 248897 292699 248931
rect 292389 248869 292437 248897
rect 292465 248869 292499 248897
rect 292527 248869 292561 248897
rect 292589 248869 292623 248897
rect 292651 248869 292699 248897
rect 292389 248835 292699 248869
rect 292389 248807 292437 248835
rect 292465 248807 292499 248835
rect 292527 248807 292561 248835
rect 292589 248807 292623 248835
rect 292651 248807 292699 248835
rect 292389 248773 292699 248807
rect 292389 248745 292437 248773
rect 292465 248745 292499 248773
rect 292527 248745 292561 248773
rect 292589 248745 292623 248773
rect 292651 248745 292699 248773
rect 292389 239959 292699 248745
rect 292389 239931 292437 239959
rect 292465 239931 292499 239959
rect 292527 239931 292561 239959
rect 292589 239931 292623 239959
rect 292651 239931 292699 239959
rect 292389 239897 292699 239931
rect 292389 239869 292437 239897
rect 292465 239869 292499 239897
rect 292527 239869 292561 239897
rect 292589 239869 292623 239897
rect 292651 239869 292699 239897
rect 292389 239835 292699 239869
rect 292389 239807 292437 239835
rect 292465 239807 292499 239835
rect 292527 239807 292561 239835
rect 292589 239807 292623 239835
rect 292651 239807 292699 239835
rect 292389 239773 292699 239807
rect 292389 239745 292437 239773
rect 292465 239745 292499 239773
rect 292527 239745 292561 239773
rect 292589 239745 292623 239773
rect 292651 239745 292699 239773
rect 292389 230959 292699 239745
rect 292389 230931 292437 230959
rect 292465 230931 292499 230959
rect 292527 230931 292561 230959
rect 292589 230931 292623 230959
rect 292651 230931 292699 230959
rect 292389 230897 292699 230931
rect 292389 230869 292437 230897
rect 292465 230869 292499 230897
rect 292527 230869 292561 230897
rect 292589 230869 292623 230897
rect 292651 230869 292699 230897
rect 292389 230835 292699 230869
rect 292389 230807 292437 230835
rect 292465 230807 292499 230835
rect 292527 230807 292561 230835
rect 292589 230807 292623 230835
rect 292651 230807 292699 230835
rect 292389 230773 292699 230807
rect 292389 230745 292437 230773
rect 292465 230745 292499 230773
rect 292527 230745 292561 230773
rect 292589 230745 292623 230773
rect 292651 230745 292699 230773
rect 292389 221959 292699 230745
rect 292389 221931 292437 221959
rect 292465 221931 292499 221959
rect 292527 221931 292561 221959
rect 292589 221931 292623 221959
rect 292651 221931 292699 221959
rect 292389 221897 292699 221931
rect 292389 221869 292437 221897
rect 292465 221869 292499 221897
rect 292527 221869 292561 221897
rect 292589 221869 292623 221897
rect 292651 221869 292699 221897
rect 292389 221835 292699 221869
rect 292389 221807 292437 221835
rect 292465 221807 292499 221835
rect 292527 221807 292561 221835
rect 292589 221807 292623 221835
rect 292651 221807 292699 221835
rect 292389 221773 292699 221807
rect 292389 221745 292437 221773
rect 292465 221745 292499 221773
rect 292527 221745 292561 221773
rect 292589 221745 292623 221773
rect 292651 221745 292699 221773
rect 292389 212959 292699 221745
rect 292389 212931 292437 212959
rect 292465 212931 292499 212959
rect 292527 212931 292561 212959
rect 292589 212931 292623 212959
rect 292651 212931 292699 212959
rect 292389 212897 292699 212931
rect 292389 212869 292437 212897
rect 292465 212869 292499 212897
rect 292527 212869 292561 212897
rect 292589 212869 292623 212897
rect 292651 212869 292699 212897
rect 292389 212835 292699 212869
rect 292389 212807 292437 212835
rect 292465 212807 292499 212835
rect 292527 212807 292561 212835
rect 292589 212807 292623 212835
rect 292651 212807 292699 212835
rect 292389 212773 292699 212807
rect 292389 212745 292437 212773
rect 292465 212745 292499 212773
rect 292527 212745 292561 212773
rect 292589 212745 292623 212773
rect 292651 212745 292699 212773
rect 292389 203959 292699 212745
rect 292389 203931 292437 203959
rect 292465 203931 292499 203959
rect 292527 203931 292561 203959
rect 292589 203931 292623 203959
rect 292651 203931 292699 203959
rect 292389 203897 292699 203931
rect 292389 203869 292437 203897
rect 292465 203869 292499 203897
rect 292527 203869 292561 203897
rect 292589 203869 292623 203897
rect 292651 203869 292699 203897
rect 292389 203835 292699 203869
rect 292389 203807 292437 203835
rect 292465 203807 292499 203835
rect 292527 203807 292561 203835
rect 292589 203807 292623 203835
rect 292651 203807 292699 203835
rect 292389 203773 292699 203807
rect 292389 203745 292437 203773
rect 292465 203745 292499 203773
rect 292527 203745 292561 203773
rect 292589 203745 292623 203773
rect 292651 203745 292699 203773
rect 292389 194959 292699 203745
rect 292389 194931 292437 194959
rect 292465 194931 292499 194959
rect 292527 194931 292561 194959
rect 292589 194931 292623 194959
rect 292651 194931 292699 194959
rect 292389 194897 292699 194931
rect 292389 194869 292437 194897
rect 292465 194869 292499 194897
rect 292527 194869 292561 194897
rect 292589 194869 292623 194897
rect 292651 194869 292699 194897
rect 292389 194835 292699 194869
rect 292389 194807 292437 194835
rect 292465 194807 292499 194835
rect 292527 194807 292561 194835
rect 292589 194807 292623 194835
rect 292651 194807 292699 194835
rect 292389 194773 292699 194807
rect 292389 194745 292437 194773
rect 292465 194745 292499 194773
rect 292527 194745 292561 194773
rect 292589 194745 292623 194773
rect 292651 194745 292699 194773
rect 292389 185959 292699 194745
rect 292389 185931 292437 185959
rect 292465 185931 292499 185959
rect 292527 185931 292561 185959
rect 292589 185931 292623 185959
rect 292651 185931 292699 185959
rect 292389 185897 292699 185931
rect 292389 185869 292437 185897
rect 292465 185869 292499 185897
rect 292527 185869 292561 185897
rect 292589 185869 292623 185897
rect 292651 185869 292699 185897
rect 292389 185835 292699 185869
rect 292389 185807 292437 185835
rect 292465 185807 292499 185835
rect 292527 185807 292561 185835
rect 292589 185807 292623 185835
rect 292651 185807 292699 185835
rect 292389 185773 292699 185807
rect 292389 185745 292437 185773
rect 292465 185745 292499 185773
rect 292527 185745 292561 185773
rect 292589 185745 292623 185773
rect 292651 185745 292699 185773
rect 292389 176959 292699 185745
rect 292389 176931 292437 176959
rect 292465 176931 292499 176959
rect 292527 176931 292561 176959
rect 292589 176931 292623 176959
rect 292651 176931 292699 176959
rect 292389 176897 292699 176931
rect 292389 176869 292437 176897
rect 292465 176869 292499 176897
rect 292527 176869 292561 176897
rect 292589 176869 292623 176897
rect 292651 176869 292699 176897
rect 292389 176835 292699 176869
rect 292389 176807 292437 176835
rect 292465 176807 292499 176835
rect 292527 176807 292561 176835
rect 292589 176807 292623 176835
rect 292651 176807 292699 176835
rect 292389 176773 292699 176807
rect 292389 176745 292437 176773
rect 292465 176745 292499 176773
rect 292527 176745 292561 176773
rect 292589 176745 292623 176773
rect 292651 176745 292699 176773
rect 292389 167959 292699 176745
rect 292389 167931 292437 167959
rect 292465 167931 292499 167959
rect 292527 167931 292561 167959
rect 292589 167931 292623 167959
rect 292651 167931 292699 167959
rect 292389 167897 292699 167931
rect 292389 167869 292437 167897
rect 292465 167869 292499 167897
rect 292527 167869 292561 167897
rect 292589 167869 292623 167897
rect 292651 167869 292699 167897
rect 292389 167835 292699 167869
rect 292389 167807 292437 167835
rect 292465 167807 292499 167835
rect 292527 167807 292561 167835
rect 292589 167807 292623 167835
rect 292651 167807 292699 167835
rect 292389 167773 292699 167807
rect 292389 167745 292437 167773
rect 292465 167745 292499 167773
rect 292527 167745 292561 167773
rect 292589 167745 292623 167773
rect 292651 167745 292699 167773
rect 292389 158959 292699 167745
rect 292389 158931 292437 158959
rect 292465 158931 292499 158959
rect 292527 158931 292561 158959
rect 292589 158931 292623 158959
rect 292651 158931 292699 158959
rect 292389 158897 292699 158931
rect 292389 158869 292437 158897
rect 292465 158869 292499 158897
rect 292527 158869 292561 158897
rect 292589 158869 292623 158897
rect 292651 158869 292699 158897
rect 292389 158835 292699 158869
rect 292389 158807 292437 158835
rect 292465 158807 292499 158835
rect 292527 158807 292561 158835
rect 292589 158807 292623 158835
rect 292651 158807 292699 158835
rect 292389 158773 292699 158807
rect 292389 158745 292437 158773
rect 292465 158745 292499 158773
rect 292527 158745 292561 158773
rect 292589 158745 292623 158773
rect 292651 158745 292699 158773
rect 292389 149959 292699 158745
rect 292389 149931 292437 149959
rect 292465 149931 292499 149959
rect 292527 149931 292561 149959
rect 292589 149931 292623 149959
rect 292651 149931 292699 149959
rect 292389 149897 292699 149931
rect 292389 149869 292437 149897
rect 292465 149869 292499 149897
rect 292527 149869 292561 149897
rect 292589 149869 292623 149897
rect 292651 149869 292699 149897
rect 292389 149835 292699 149869
rect 292389 149807 292437 149835
rect 292465 149807 292499 149835
rect 292527 149807 292561 149835
rect 292589 149807 292623 149835
rect 292651 149807 292699 149835
rect 292389 149773 292699 149807
rect 292389 149745 292437 149773
rect 292465 149745 292499 149773
rect 292527 149745 292561 149773
rect 292589 149745 292623 149773
rect 292651 149745 292699 149773
rect 292389 140959 292699 149745
rect 292389 140931 292437 140959
rect 292465 140931 292499 140959
rect 292527 140931 292561 140959
rect 292589 140931 292623 140959
rect 292651 140931 292699 140959
rect 292389 140897 292699 140931
rect 292389 140869 292437 140897
rect 292465 140869 292499 140897
rect 292527 140869 292561 140897
rect 292589 140869 292623 140897
rect 292651 140869 292699 140897
rect 292389 140835 292699 140869
rect 292389 140807 292437 140835
rect 292465 140807 292499 140835
rect 292527 140807 292561 140835
rect 292589 140807 292623 140835
rect 292651 140807 292699 140835
rect 292389 140773 292699 140807
rect 292389 140745 292437 140773
rect 292465 140745 292499 140773
rect 292527 140745 292561 140773
rect 292589 140745 292623 140773
rect 292651 140745 292699 140773
rect 292389 131959 292699 140745
rect 292389 131931 292437 131959
rect 292465 131931 292499 131959
rect 292527 131931 292561 131959
rect 292589 131931 292623 131959
rect 292651 131931 292699 131959
rect 292389 131897 292699 131931
rect 292389 131869 292437 131897
rect 292465 131869 292499 131897
rect 292527 131869 292561 131897
rect 292589 131869 292623 131897
rect 292651 131869 292699 131897
rect 292389 131835 292699 131869
rect 292389 131807 292437 131835
rect 292465 131807 292499 131835
rect 292527 131807 292561 131835
rect 292589 131807 292623 131835
rect 292651 131807 292699 131835
rect 292389 131773 292699 131807
rect 292389 131745 292437 131773
rect 292465 131745 292499 131773
rect 292527 131745 292561 131773
rect 292589 131745 292623 131773
rect 292651 131745 292699 131773
rect 292389 122959 292699 131745
rect 292389 122931 292437 122959
rect 292465 122931 292499 122959
rect 292527 122931 292561 122959
rect 292589 122931 292623 122959
rect 292651 122931 292699 122959
rect 292389 122897 292699 122931
rect 292389 122869 292437 122897
rect 292465 122869 292499 122897
rect 292527 122869 292561 122897
rect 292589 122869 292623 122897
rect 292651 122869 292699 122897
rect 292389 122835 292699 122869
rect 292389 122807 292437 122835
rect 292465 122807 292499 122835
rect 292527 122807 292561 122835
rect 292589 122807 292623 122835
rect 292651 122807 292699 122835
rect 292389 122773 292699 122807
rect 292389 122745 292437 122773
rect 292465 122745 292499 122773
rect 292527 122745 292561 122773
rect 292589 122745 292623 122773
rect 292651 122745 292699 122773
rect 292389 113959 292699 122745
rect 292389 113931 292437 113959
rect 292465 113931 292499 113959
rect 292527 113931 292561 113959
rect 292589 113931 292623 113959
rect 292651 113931 292699 113959
rect 292389 113897 292699 113931
rect 292389 113869 292437 113897
rect 292465 113869 292499 113897
rect 292527 113869 292561 113897
rect 292589 113869 292623 113897
rect 292651 113869 292699 113897
rect 292389 113835 292699 113869
rect 292389 113807 292437 113835
rect 292465 113807 292499 113835
rect 292527 113807 292561 113835
rect 292589 113807 292623 113835
rect 292651 113807 292699 113835
rect 292389 113773 292699 113807
rect 292389 113745 292437 113773
rect 292465 113745 292499 113773
rect 292527 113745 292561 113773
rect 292589 113745 292623 113773
rect 292651 113745 292699 113773
rect 292389 104959 292699 113745
rect 292389 104931 292437 104959
rect 292465 104931 292499 104959
rect 292527 104931 292561 104959
rect 292589 104931 292623 104959
rect 292651 104931 292699 104959
rect 292389 104897 292699 104931
rect 292389 104869 292437 104897
rect 292465 104869 292499 104897
rect 292527 104869 292561 104897
rect 292589 104869 292623 104897
rect 292651 104869 292699 104897
rect 292389 104835 292699 104869
rect 292389 104807 292437 104835
rect 292465 104807 292499 104835
rect 292527 104807 292561 104835
rect 292589 104807 292623 104835
rect 292651 104807 292699 104835
rect 292389 104773 292699 104807
rect 292389 104745 292437 104773
rect 292465 104745 292499 104773
rect 292527 104745 292561 104773
rect 292589 104745 292623 104773
rect 292651 104745 292699 104773
rect 292389 95959 292699 104745
rect 292389 95931 292437 95959
rect 292465 95931 292499 95959
rect 292527 95931 292561 95959
rect 292589 95931 292623 95959
rect 292651 95931 292699 95959
rect 292389 95897 292699 95931
rect 292389 95869 292437 95897
rect 292465 95869 292499 95897
rect 292527 95869 292561 95897
rect 292589 95869 292623 95897
rect 292651 95869 292699 95897
rect 292389 95835 292699 95869
rect 292389 95807 292437 95835
rect 292465 95807 292499 95835
rect 292527 95807 292561 95835
rect 292589 95807 292623 95835
rect 292651 95807 292699 95835
rect 292389 95773 292699 95807
rect 292389 95745 292437 95773
rect 292465 95745 292499 95773
rect 292527 95745 292561 95773
rect 292589 95745 292623 95773
rect 292651 95745 292699 95773
rect 292389 86959 292699 95745
rect 292389 86931 292437 86959
rect 292465 86931 292499 86959
rect 292527 86931 292561 86959
rect 292589 86931 292623 86959
rect 292651 86931 292699 86959
rect 292389 86897 292699 86931
rect 292389 86869 292437 86897
rect 292465 86869 292499 86897
rect 292527 86869 292561 86897
rect 292589 86869 292623 86897
rect 292651 86869 292699 86897
rect 292389 86835 292699 86869
rect 292389 86807 292437 86835
rect 292465 86807 292499 86835
rect 292527 86807 292561 86835
rect 292589 86807 292623 86835
rect 292651 86807 292699 86835
rect 292389 86773 292699 86807
rect 292389 86745 292437 86773
rect 292465 86745 292499 86773
rect 292527 86745 292561 86773
rect 292589 86745 292623 86773
rect 292651 86745 292699 86773
rect 292389 77959 292699 86745
rect 292389 77931 292437 77959
rect 292465 77931 292499 77959
rect 292527 77931 292561 77959
rect 292589 77931 292623 77959
rect 292651 77931 292699 77959
rect 292389 77897 292699 77931
rect 292389 77869 292437 77897
rect 292465 77869 292499 77897
rect 292527 77869 292561 77897
rect 292589 77869 292623 77897
rect 292651 77869 292699 77897
rect 292389 77835 292699 77869
rect 292389 77807 292437 77835
rect 292465 77807 292499 77835
rect 292527 77807 292561 77835
rect 292589 77807 292623 77835
rect 292651 77807 292699 77835
rect 292389 77773 292699 77807
rect 292389 77745 292437 77773
rect 292465 77745 292499 77773
rect 292527 77745 292561 77773
rect 292589 77745 292623 77773
rect 292651 77745 292699 77773
rect 292389 68959 292699 77745
rect 292389 68931 292437 68959
rect 292465 68931 292499 68959
rect 292527 68931 292561 68959
rect 292589 68931 292623 68959
rect 292651 68931 292699 68959
rect 292389 68897 292699 68931
rect 292389 68869 292437 68897
rect 292465 68869 292499 68897
rect 292527 68869 292561 68897
rect 292589 68869 292623 68897
rect 292651 68869 292699 68897
rect 292389 68835 292699 68869
rect 292389 68807 292437 68835
rect 292465 68807 292499 68835
rect 292527 68807 292561 68835
rect 292589 68807 292623 68835
rect 292651 68807 292699 68835
rect 292389 68773 292699 68807
rect 292389 68745 292437 68773
rect 292465 68745 292499 68773
rect 292527 68745 292561 68773
rect 292589 68745 292623 68773
rect 292651 68745 292699 68773
rect 292389 59959 292699 68745
rect 292389 59931 292437 59959
rect 292465 59931 292499 59959
rect 292527 59931 292561 59959
rect 292589 59931 292623 59959
rect 292651 59931 292699 59959
rect 292389 59897 292699 59931
rect 292389 59869 292437 59897
rect 292465 59869 292499 59897
rect 292527 59869 292561 59897
rect 292589 59869 292623 59897
rect 292651 59869 292699 59897
rect 292389 59835 292699 59869
rect 292389 59807 292437 59835
rect 292465 59807 292499 59835
rect 292527 59807 292561 59835
rect 292589 59807 292623 59835
rect 292651 59807 292699 59835
rect 292389 59773 292699 59807
rect 292389 59745 292437 59773
rect 292465 59745 292499 59773
rect 292527 59745 292561 59773
rect 292589 59745 292623 59773
rect 292651 59745 292699 59773
rect 292389 50959 292699 59745
rect 292389 50931 292437 50959
rect 292465 50931 292499 50959
rect 292527 50931 292561 50959
rect 292589 50931 292623 50959
rect 292651 50931 292699 50959
rect 292389 50897 292699 50931
rect 292389 50869 292437 50897
rect 292465 50869 292499 50897
rect 292527 50869 292561 50897
rect 292589 50869 292623 50897
rect 292651 50869 292699 50897
rect 292389 50835 292699 50869
rect 292389 50807 292437 50835
rect 292465 50807 292499 50835
rect 292527 50807 292561 50835
rect 292589 50807 292623 50835
rect 292651 50807 292699 50835
rect 292389 50773 292699 50807
rect 292389 50745 292437 50773
rect 292465 50745 292499 50773
rect 292527 50745 292561 50773
rect 292589 50745 292623 50773
rect 292651 50745 292699 50773
rect 292389 41959 292699 50745
rect 292389 41931 292437 41959
rect 292465 41931 292499 41959
rect 292527 41931 292561 41959
rect 292589 41931 292623 41959
rect 292651 41931 292699 41959
rect 292389 41897 292699 41931
rect 292389 41869 292437 41897
rect 292465 41869 292499 41897
rect 292527 41869 292561 41897
rect 292589 41869 292623 41897
rect 292651 41869 292699 41897
rect 292389 41835 292699 41869
rect 292389 41807 292437 41835
rect 292465 41807 292499 41835
rect 292527 41807 292561 41835
rect 292589 41807 292623 41835
rect 292651 41807 292699 41835
rect 292389 41773 292699 41807
rect 292389 41745 292437 41773
rect 292465 41745 292499 41773
rect 292527 41745 292561 41773
rect 292589 41745 292623 41773
rect 292651 41745 292699 41773
rect 292389 32959 292699 41745
rect 292389 32931 292437 32959
rect 292465 32931 292499 32959
rect 292527 32931 292561 32959
rect 292589 32931 292623 32959
rect 292651 32931 292699 32959
rect 292389 32897 292699 32931
rect 292389 32869 292437 32897
rect 292465 32869 292499 32897
rect 292527 32869 292561 32897
rect 292589 32869 292623 32897
rect 292651 32869 292699 32897
rect 292389 32835 292699 32869
rect 292389 32807 292437 32835
rect 292465 32807 292499 32835
rect 292527 32807 292561 32835
rect 292589 32807 292623 32835
rect 292651 32807 292699 32835
rect 292389 32773 292699 32807
rect 292389 32745 292437 32773
rect 292465 32745 292499 32773
rect 292527 32745 292561 32773
rect 292589 32745 292623 32773
rect 292651 32745 292699 32773
rect 292389 23959 292699 32745
rect 292389 23931 292437 23959
rect 292465 23931 292499 23959
rect 292527 23931 292561 23959
rect 292589 23931 292623 23959
rect 292651 23931 292699 23959
rect 292389 23897 292699 23931
rect 292389 23869 292437 23897
rect 292465 23869 292499 23897
rect 292527 23869 292561 23897
rect 292589 23869 292623 23897
rect 292651 23869 292699 23897
rect 292389 23835 292699 23869
rect 292389 23807 292437 23835
rect 292465 23807 292499 23835
rect 292527 23807 292561 23835
rect 292589 23807 292623 23835
rect 292651 23807 292699 23835
rect 292389 23773 292699 23807
rect 292389 23745 292437 23773
rect 292465 23745 292499 23773
rect 292527 23745 292561 23773
rect 292589 23745 292623 23773
rect 292651 23745 292699 23773
rect 292389 14959 292699 23745
rect 292389 14931 292437 14959
rect 292465 14931 292499 14959
rect 292527 14931 292561 14959
rect 292589 14931 292623 14959
rect 292651 14931 292699 14959
rect 292389 14897 292699 14931
rect 292389 14869 292437 14897
rect 292465 14869 292499 14897
rect 292527 14869 292561 14897
rect 292589 14869 292623 14897
rect 292651 14869 292699 14897
rect 292389 14835 292699 14869
rect 292389 14807 292437 14835
rect 292465 14807 292499 14835
rect 292527 14807 292561 14835
rect 292589 14807 292623 14835
rect 292651 14807 292699 14835
rect 292389 14773 292699 14807
rect 292389 14745 292437 14773
rect 292465 14745 292499 14773
rect 292527 14745 292561 14773
rect 292589 14745 292623 14773
rect 292651 14745 292699 14773
rect 292389 5959 292699 14745
rect 292389 5931 292437 5959
rect 292465 5931 292499 5959
rect 292527 5931 292561 5959
rect 292589 5931 292623 5959
rect 292651 5931 292699 5959
rect 292389 5897 292699 5931
rect 292389 5869 292437 5897
rect 292465 5869 292499 5897
rect 292527 5869 292561 5897
rect 292589 5869 292623 5897
rect 292651 5869 292699 5897
rect 292389 5835 292699 5869
rect 292389 5807 292437 5835
rect 292465 5807 292499 5835
rect 292527 5807 292561 5835
rect 292589 5807 292623 5835
rect 292651 5807 292699 5835
rect 292389 5773 292699 5807
rect 292389 5745 292437 5773
rect 292465 5745 292499 5773
rect 292527 5745 292561 5773
rect 292589 5745 292623 5773
rect 292651 5745 292699 5773
rect 292389 424 292699 5745
rect 299208 299190 299518 299238
rect 299208 299162 299256 299190
rect 299284 299162 299318 299190
rect 299346 299162 299380 299190
rect 299408 299162 299442 299190
rect 299470 299162 299518 299190
rect 299208 299128 299518 299162
rect 299208 299100 299256 299128
rect 299284 299100 299318 299128
rect 299346 299100 299380 299128
rect 299408 299100 299442 299128
rect 299470 299100 299518 299128
rect 299208 299066 299518 299100
rect 299208 299038 299256 299066
rect 299284 299038 299318 299066
rect 299346 299038 299380 299066
rect 299408 299038 299442 299066
rect 299470 299038 299518 299066
rect 299208 299004 299518 299038
rect 299208 298976 299256 299004
rect 299284 298976 299318 299004
rect 299346 298976 299380 299004
rect 299408 298976 299442 299004
rect 299470 298976 299518 299004
rect 299208 290959 299518 298976
rect 299208 290931 299256 290959
rect 299284 290931 299318 290959
rect 299346 290931 299380 290959
rect 299408 290931 299442 290959
rect 299470 290931 299518 290959
rect 299208 290897 299518 290931
rect 299208 290869 299256 290897
rect 299284 290869 299318 290897
rect 299346 290869 299380 290897
rect 299408 290869 299442 290897
rect 299470 290869 299518 290897
rect 299208 290835 299518 290869
rect 299208 290807 299256 290835
rect 299284 290807 299318 290835
rect 299346 290807 299380 290835
rect 299408 290807 299442 290835
rect 299470 290807 299518 290835
rect 299208 290773 299518 290807
rect 299208 290745 299256 290773
rect 299284 290745 299318 290773
rect 299346 290745 299380 290773
rect 299408 290745 299442 290773
rect 299470 290745 299518 290773
rect 299208 281959 299518 290745
rect 299208 281931 299256 281959
rect 299284 281931 299318 281959
rect 299346 281931 299380 281959
rect 299408 281931 299442 281959
rect 299470 281931 299518 281959
rect 299208 281897 299518 281931
rect 299208 281869 299256 281897
rect 299284 281869 299318 281897
rect 299346 281869 299380 281897
rect 299408 281869 299442 281897
rect 299470 281869 299518 281897
rect 299208 281835 299518 281869
rect 299208 281807 299256 281835
rect 299284 281807 299318 281835
rect 299346 281807 299380 281835
rect 299408 281807 299442 281835
rect 299470 281807 299518 281835
rect 299208 281773 299518 281807
rect 299208 281745 299256 281773
rect 299284 281745 299318 281773
rect 299346 281745 299380 281773
rect 299408 281745 299442 281773
rect 299470 281745 299518 281773
rect 299208 272959 299518 281745
rect 299208 272931 299256 272959
rect 299284 272931 299318 272959
rect 299346 272931 299380 272959
rect 299408 272931 299442 272959
rect 299470 272931 299518 272959
rect 299208 272897 299518 272931
rect 299208 272869 299256 272897
rect 299284 272869 299318 272897
rect 299346 272869 299380 272897
rect 299408 272869 299442 272897
rect 299470 272869 299518 272897
rect 299208 272835 299518 272869
rect 299208 272807 299256 272835
rect 299284 272807 299318 272835
rect 299346 272807 299380 272835
rect 299408 272807 299442 272835
rect 299470 272807 299518 272835
rect 299208 272773 299518 272807
rect 299208 272745 299256 272773
rect 299284 272745 299318 272773
rect 299346 272745 299380 272773
rect 299408 272745 299442 272773
rect 299470 272745 299518 272773
rect 299208 263959 299518 272745
rect 299208 263931 299256 263959
rect 299284 263931 299318 263959
rect 299346 263931 299380 263959
rect 299408 263931 299442 263959
rect 299470 263931 299518 263959
rect 299208 263897 299518 263931
rect 299208 263869 299256 263897
rect 299284 263869 299318 263897
rect 299346 263869 299380 263897
rect 299408 263869 299442 263897
rect 299470 263869 299518 263897
rect 299208 263835 299518 263869
rect 299208 263807 299256 263835
rect 299284 263807 299318 263835
rect 299346 263807 299380 263835
rect 299408 263807 299442 263835
rect 299470 263807 299518 263835
rect 299208 263773 299518 263807
rect 299208 263745 299256 263773
rect 299284 263745 299318 263773
rect 299346 263745 299380 263773
rect 299408 263745 299442 263773
rect 299470 263745 299518 263773
rect 299208 254959 299518 263745
rect 299208 254931 299256 254959
rect 299284 254931 299318 254959
rect 299346 254931 299380 254959
rect 299408 254931 299442 254959
rect 299470 254931 299518 254959
rect 299208 254897 299518 254931
rect 299208 254869 299256 254897
rect 299284 254869 299318 254897
rect 299346 254869 299380 254897
rect 299408 254869 299442 254897
rect 299470 254869 299518 254897
rect 299208 254835 299518 254869
rect 299208 254807 299256 254835
rect 299284 254807 299318 254835
rect 299346 254807 299380 254835
rect 299408 254807 299442 254835
rect 299470 254807 299518 254835
rect 299208 254773 299518 254807
rect 299208 254745 299256 254773
rect 299284 254745 299318 254773
rect 299346 254745 299380 254773
rect 299408 254745 299442 254773
rect 299470 254745 299518 254773
rect 299208 245959 299518 254745
rect 299208 245931 299256 245959
rect 299284 245931 299318 245959
rect 299346 245931 299380 245959
rect 299408 245931 299442 245959
rect 299470 245931 299518 245959
rect 299208 245897 299518 245931
rect 299208 245869 299256 245897
rect 299284 245869 299318 245897
rect 299346 245869 299380 245897
rect 299408 245869 299442 245897
rect 299470 245869 299518 245897
rect 299208 245835 299518 245869
rect 299208 245807 299256 245835
rect 299284 245807 299318 245835
rect 299346 245807 299380 245835
rect 299408 245807 299442 245835
rect 299470 245807 299518 245835
rect 299208 245773 299518 245807
rect 299208 245745 299256 245773
rect 299284 245745 299318 245773
rect 299346 245745 299380 245773
rect 299408 245745 299442 245773
rect 299470 245745 299518 245773
rect 299208 236959 299518 245745
rect 299208 236931 299256 236959
rect 299284 236931 299318 236959
rect 299346 236931 299380 236959
rect 299408 236931 299442 236959
rect 299470 236931 299518 236959
rect 299208 236897 299518 236931
rect 299208 236869 299256 236897
rect 299284 236869 299318 236897
rect 299346 236869 299380 236897
rect 299408 236869 299442 236897
rect 299470 236869 299518 236897
rect 299208 236835 299518 236869
rect 299208 236807 299256 236835
rect 299284 236807 299318 236835
rect 299346 236807 299380 236835
rect 299408 236807 299442 236835
rect 299470 236807 299518 236835
rect 299208 236773 299518 236807
rect 299208 236745 299256 236773
rect 299284 236745 299318 236773
rect 299346 236745 299380 236773
rect 299408 236745 299442 236773
rect 299470 236745 299518 236773
rect 299208 227959 299518 236745
rect 299208 227931 299256 227959
rect 299284 227931 299318 227959
rect 299346 227931 299380 227959
rect 299408 227931 299442 227959
rect 299470 227931 299518 227959
rect 299208 227897 299518 227931
rect 299208 227869 299256 227897
rect 299284 227869 299318 227897
rect 299346 227869 299380 227897
rect 299408 227869 299442 227897
rect 299470 227869 299518 227897
rect 299208 227835 299518 227869
rect 299208 227807 299256 227835
rect 299284 227807 299318 227835
rect 299346 227807 299380 227835
rect 299408 227807 299442 227835
rect 299470 227807 299518 227835
rect 299208 227773 299518 227807
rect 299208 227745 299256 227773
rect 299284 227745 299318 227773
rect 299346 227745 299380 227773
rect 299408 227745 299442 227773
rect 299470 227745 299518 227773
rect 299208 218959 299518 227745
rect 299208 218931 299256 218959
rect 299284 218931 299318 218959
rect 299346 218931 299380 218959
rect 299408 218931 299442 218959
rect 299470 218931 299518 218959
rect 299208 218897 299518 218931
rect 299208 218869 299256 218897
rect 299284 218869 299318 218897
rect 299346 218869 299380 218897
rect 299408 218869 299442 218897
rect 299470 218869 299518 218897
rect 299208 218835 299518 218869
rect 299208 218807 299256 218835
rect 299284 218807 299318 218835
rect 299346 218807 299380 218835
rect 299408 218807 299442 218835
rect 299470 218807 299518 218835
rect 299208 218773 299518 218807
rect 299208 218745 299256 218773
rect 299284 218745 299318 218773
rect 299346 218745 299380 218773
rect 299408 218745 299442 218773
rect 299470 218745 299518 218773
rect 299208 209959 299518 218745
rect 299208 209931 299256 209959
rect 299284 209931 299318 209959
rect 299346 209931 299380 209959
rect 299408 209931 299442 209959
rect 299470 209931 299518 209959
rect 299208 209897 299518 209931
rect 299208 209869 299256 209897
rect 299284 209869 299318 209897
rect 299346 209869 299380 209897
rect 299408 209869 299442 209897
rect 299470 209869 299518 209897
rect 299208 209835 299518 209869
rect 299208 209807 299256 209835
rect 299284 209807 299318 209835
rect 299346 209807 299380 209835
rect 299408 209807 299442 209835
rect 299470 209807 299518 209835
rect 299208 209773 299518 209807
rect 299208 209745 299256 209773
rect 299284 209745 299318 209773
rect 299346 209745 299380 209773
rect 299408 209745 299442 209773
rect 299470 209745 299518 209773
rect 299208 200959 299518 209745
rect 299208 200931 299256 200959
rect 299284 200931 299318 200959
rect 299346 200931 299380 200959
rect 299408 200931 299442 200959
rect 299470 200931 299518 200959
rect 299208 200897 299518 200931
rect 299208 200869 299256 200897
rect 299284 200869 299318 200897
rect 299346 200869 299380 200897
rect 299408 200869 299442 200897
rect 299470 200869 299518 200897
rect 299208 200835 299518 200869
rect 299208 200807 299256 200835
rect 299284 200807 299318 200835
rect 299346 200807 299380 200835
rect 299408 200807 299442 200835
rect 299470 200807 299518 200835
rect 299208 200773 299518 200807
rect 299208 200745 299256 200773
rect 299284 200745 299318 200773
rect 299346 200745 299380 200773
rect 299408 200745 299442 200773
rect 299470 200745 299518 200773
rect 299208 191959 299518 200745
rect 299208 191931 299256 191959
rect 299284 191931 299318 191959
rect 299346 191931 299380 191959
rect 299408 191931 299442 191959
rect 299470 191931 299518 191959
rect 299208 191897 299518 191931
rect 299208 191869 299256 191897
rect 299284 191869 299318 191897
rect 299346 191869 299380 191897
rect 299408 191869 299442 191897
rect 299470 191869 299518 191897
rect 299208 191835 299518 191869
rect 299208 191807 299256 191835
rect 299284 191807 299318 191835
rect 299346 191807 299380 191835
rect 299408 191807 299442 191835
rect 299470 191807 299518 191835
rect 299208 191773 299518 191807
rect 299208 191745 299256 191773
rect 299284 191745 299318 191773
rect 299346 191745 299380 191773
rect 299408 191745 299442 191773
rect 299470 191745 299518 191773
rect 299208 182959 299518 191745
rect 299208 182931 299256 182959
rect 299284 182931 299318 182959
rect 299346 182931 299380 182959
rect 299408 182931 299442 182959
rect 299470 182931 299518 182959
rect 299208 182897 299518 182931
rect 299208 182869 299256 182897
rect 299284 182869 299318 182897
rect 299346 182869 299380 182897
rect 299408 182869 299442 182897
rect 299470 182869 299518 182897
rect 299208 182835 299518 182869
rect 299208 182807 299256 182835
rect 299284 182807 299318 182835
rect 299346 182807 299380 182835
rect 299408 182807 299442 182835
rect 299470 182807 299518 182835
rect 299208 182773 299518 182807
rect 299208 182745 299256 182773
rect 299284 182745 299318 182773
rect 299346 182745 299380 182773
rect 299408 182745 299442 182773
rect 299470 182745 299518 182773
rect 299208 173959 299518 182745
rect 299208 173931 299256 173959
rect 299284 173931 299318 173959
rect 299346 173931 299380 173959
rect 299408 173931 299442 173959
rect 299470 173931 299518 173959
rect 299208 173897 299518 173931
rect 299208 173869 299256 173897
rect 299284 173869 299318 173897
rect 299346 173869 299380 173897
rect 299408 173869 299442 173897
rect 299470 173869 299518 173897
rect 299208 173835 299518 173869
rect 299208 173807 299256 173835
rect 299284 173807 299318 173835
rect 299346 173807 299380 173835
rect 299408 173807 299442 173835
rect 299470 173807 299518 173835
rect 299208 173773 299518 173807
rect 299208 173745 299256 173773
rect 299284 173745 299318 173773
rect 299346 173745 299380 173773
rect 299408 173745 299442 173773
rect 299470 173745 299518 173773
rect 299208 164959 299518 173745
rect 299208 164931 299256 164959
rect 299284 164931 299318 164959
rect 299346 164931 299380 164959
rect 299408 164931 299442 164959
rect 299470 164931 299518 164959
rect 299208 164897 299518 164931
rect 299208 164869 299256 164897
rect 299284 164869 299318 164897
rect 299346 164869 299380 164897
rect 299408 164869 299442 164897
rect 299470 164869 299518 164897
rect 299208 164835 299518 164869
rect 299208 164807 299256 164835
rect 299284 164807 299318 164835
rect 299346 164807 299380 164835
rect 299408 164807 299442 164835
rect 299470 164807 299518 164835
rect 299208 164773 299518 164807
rect 299208 164745 299256 164773
rect 299284 164745 299318 164773
rect 299346 164745 299380 164773
rect 299408 164745 299442 164773
rect 299470 164745 299518 164773
rect 299208 155959 299518 164745
rect 299208 155931 299256 155959
rect 299284 155931 299318 155959
rect 299346 155931 299380 155959
rect 299408 155931 299442 155959
rect 299470 155931 299518 155959
rect 299208 155897 299518 155931
rect 299208 155869 299256 155897
rect 299284 155869 299318 155897
rect 299346 155869 299380 155897
rect 299408 155869 299442 155897
rect 299470 155869 299518 155897
rect 299208 155835 299518 155869
rect 299208 155807 299256 155835
rect 299284 155807 299318 155835
rect 299346 155807 299380 155835
rect 299408 155807 299442 155835
rect 299470 155807 299518 155835
rect 299208 155773 299518 155807
rect 299208 155745 299256 155773
rect 299284 155745 299318 155773
rect 299346 155745 299380 155773
rect 299408 155745 299442 155773
rect 299470 155745 299518 155773
rect 299208 146959 299518 155745
rect 299208 146931 299256 146959
rect 299284 146931 299318 146959
rect 299346 146931 299380 146959
rect 299408 146931 299442 146959
rect 299470 146931 299518 146959
rect 299208 146897 299518 146931
rect 299208 146869 299256 146897
rect 299284 146869 299318 146897
rect 299346 146869 299380 146897
rect 299408 146869 299442 146897
rect 299470 146869 299518 146897
rect 299208 146835 299518 146869
rect 299208 146807 299256 146835
rect 299284 146807 299318 146835
rect 299346 146807 299380 146835
rect 299408 146807 299442 146835
rect 299470 146807 299518 146835
rect 299208 146773 299518 146807
rect 299208 146745 299256 146773
rect 299284 146745 299318 146773
rect 299346 146745 299380 146773
rect 299408 146745 299442 146773
rect 299470 146745 299518 146773
rect 299208 137959 299518 146745
rect 299208 137931 299256 137959
rect 299284 137931 299318 137959
rect 299346 137931 299380 137959
rect 299408 137931 299442 137959
rect 299470 137931 299518 137959
rect 299208 137897 299518 137931
rect 299208 137869 299256 137897
rect 299284 137869 299318 137897
rect 299346 137869 299380 137897
rect 299408 137869 299442 137897
rect 299470 137869 299518 137897
rect 299208 137835 299518 137869
rect 299208 137807 299256 137835
rect 299284 137807 299318 137835
rect 299346 137807 299380 137835
rect 299408 137807 299442 137835
rect 299470 137807 299518 137835
rect 299208 137773 299518 137807
rect 299208 137745 299256 137773
rect 299284 137745 299318 137773
rect 299346 137745 299380 137773
rect 299408 137745 299442 137773
rect 299470 137745 299518 137773
rect 299208 128959 299518 137745
rect 299208 128931 299256 128959
rect 299284 128931 299318 128959
rect 299346 128931 299380 128959
rect 299408 128931 299442 128959
rect 299470 128931 299518 128959
rect 299208 128897 299518 128931
rect 299208 128869 299256 128897
rect 299284 128869 299318 128897
rect 299346 128869 299380 128897
rect 299408 128869 299442 128897
rect 299470 128869 299518 128897
rect 299208 128835 299518 128869
rect 299208 128807 299256 128835
rect 299284 128807 299318 128835
rect 299346 128807 299380 128835
rect 299408 128807 299442 128835
rect 299470 128807 299518 128835
rect 299208 128773 299518 128807
rect 299208 128745 299256 128773
rect 299284 128745 299318 128773
rect 299346 128745 299380 128773
rect 299408 128745 299442 128773
rect 299470 128745 299518 128773
rect 299208 119959 299518 128745
rect 299208 119931 299256 119959
rect 299284 119931 299318 119959
rect 299346 119931 299380 119959
rect 299408 119931 299442 119959
rect 299470 119931 299518 119959
rect 299208 119897 299518 119931
rect 299208 119869 299256 119897
rect 299284 119869 299318 119897
rect 299346 119869 299380 119897
rect 299408 119869 299442 119897
rect 299470 119869 299518 119897
rect 299208 119835 299518 119869
rect 299208 119807 299256 119835
rect 299284 119807 299318 119835
rect 299346 119807 299380 119835
rect 299408 119807 299442 119835
rect 299470 119807 299518 119835
rect 299208 119773 299518 119807
rect 299208 119745 299256 119773
rect 299284 119745 299318 119773
rect 299346 119745 299380 119773
rect 299408 119745 299442 119773
rect 299470 119745 299518 119773
rect 299208 110959 299518 119745
rect 299208 110931 299256 110959
rect 299284 110931 299318 110959
rect 299346 110931 299380 110959
rect 299408 110931 299442 110959
rect 299470 110931 299518 110959
rect 299208 110897 299518 110931
rect 299208 110869 299256 110897
rect 299284 110869 299318 110897
rect 299346 110869 299380 110897
rect 299408 110869 299442 110897
rect 299470 110869 299518 110897
rect 299208 110835 299518 110869
rect 299208 110807 299256 110835
rect 299284 110807 299318 110835
rect 299346 110807 299380 110835
rect 299408 110807 299442 110835
rect 299470 110807 299518 110835
rect 299208 110773 299518 110807
rect 299208 110745 299256 110773
rect 299284 110745 299318 110773
rect 299346 110745 299380 110773
rect 299408 110745 299442 110773
rect 299470 110745 299518 110773
rect 299208 101959 299518 110745
rect 299208 101931 299256 101959
rect 299284 101931 299318 101959
rect 299346 101931 299380 101959
rect 299408 101931 299442 101959
rect 299470 101931 299518 101959
rect 299208 101897 299518 101931
rect 299208 101869 299256 101897
rect 299284 101869 299318 101897
rect 299346 101869 299380 101897
rect 299408 101869 299442 101897
rect 299470 101869 299518 101897
rect 299208 101835 299518 101869
rect 299208 101807 299256 101835
rect 299284 101807 299318 101835
rect 299346 101807 299380 101835
rect 299408 101807 299442 101835
rect 299470 101807 299518 101835
rect 299208 101773 299518 101807
rect 299208 101745 299256 101773
rect 299284 101745 299318 101773
rect 299346 101745 299380 101773
rect 299408 101745 299442 101773
rect 299470 101745 299518 101773
rect 299208 92959 299518 101745
rect 299208 92931 299256 92959
rect 299284 92931 299318 92959
rect 299346 92931 299380 92959
rect 299408 92931 299442 92959
rect 299470 92931 299518 92959
rect 299208 92897 299518 92931
rect 299208 92869 299256 92897
rect 299284 92869 299318 92897
rect 299346 92869 299380 92897
rect 299408 92869 299442 92897
rect 299470 92869 299518 92897
rect 299208 92835 299518 92869
rect 299208 92807 299256 92835
rect 299284 92807 299318 92835
rect 299346 92807 299380 92835
rect 299408 92807 299442 92835
rect 299470 92807 299518 92835
rect 299208 92773 299518 92807
rect 299208 92745 299256 92773
rect 299284 92745 299318 92773
rect 299346 92745 299380 92773
rect 299408 92745 299442 92773
rect 299470 92745 299518 92773
rect 299208 83959 299518 92745
rect 299208 83931 299256 83959
rect 299284 83931 299318 83959
rect 299346 83931 299380 83959
rect 299408 83931 299442 83959
rect 299470 83931 299518 83959
rect 299208 83897 299518 83931
rect 299208 83869 299256 83897
rect 299284 83869 299318 83897
rect 299346 83869 299380 83897
rect 299408 83869 299442 83897
rect 299470 83869 299518 83897
rect 299208 83835 299518 83869
rect 299208 83807 299256 83835
rect 299284 83807 299318 83835
rect 299346 83807 299380 83835
rect 299408 83807 299442 83835
rect 299470 83807 299518 83835
rect 299208 83773 299518 83807
rect 299208 83745 299256 83773
rect 299284 83745 299318 83773
rect 299346 83745 299380 83773
rect 299408 83745 299442 83773
rect 299470 83745 299518 83773
rect 299208 74959 299518 83745
rect 299208 74931 299256 74959
rect 299284 74931 299318 74959
rect 299346 74931 299380 74959
rect 299408 74931 299442 74959
rect 299470 74931 299518 74959
rect 299208 74897 299518 74931
rect 299208 74869 299256 74897
rect 299284 74869 299318 74897
rect 299346 74869 299380 74897
rect 299408 74869 299442 74897
rect 299470 74869 299518 74897
rect 299208 74835 299518 74869
rect 299208 74807 299256 74835
rect 299284 74807 299318 74835
rect 299346 74807 299380 74835
rect 299408 74807 299442 74835
rect 299470 74807 299518 74835
rect 299208 74773 299518 74807
rect 299208 74745 299256 74773
rect 299284 74745 299318 74773
rect 299346 74745 299380 74773
rect 299408 74745 299442 74773
rect 299470 74745 299518 74773
rect 299208 65959 299518 74745
rect 299208 65931 299256 65959
rect 299284 65931 299318 65959
rect 299346 65931 299380 65959
rect 299408 65931 299442 65959
rect 299470 65931 299518 65959
rect 299208 65897 299518 65931
rect 299208 65869 299256 65897
rect 299284 65869 299318 65897
rect 299346 65869 299380 65897
rect 299408 65869 299442 65897
rect 299470 65869 299518 65897
rect 299208 65835 299518 65869
rect 299208 65807 299256 65835
rect 299284 65807 299318 65835
rect 299346 65807 299380 65835
rect 299408 65807 299442 65835
rect 299470 65807 299518 65835
rect 299208 65773 299518 65807
rect 299208 65745 299256 65773
rect 299284 65745 299318 65773
rect 299346 65745 299380 65773
rect 299408 65745 299442 65773
rect 299470 65745 299518 65773
rect 299208 56959 299518 65745
rect 299208 56931 299256 56959
rect 299284 56931 299318 56959
rect 299346 56931 299380 56959
rect 299408 56931 299442 56959
rect 299470 56931 299518 56959
rect 299208 56897 299518 56931
rect 299208 56869 299256 56897
rect 299284 56869 299318 56897
rect 299346 56869 299380 56897
rect 299408 56869 299442 56897
rect 299470 56869 299518 56897
rect 299208 56835 299518 56869
rect 299208 56807 299256 56835
rect 299284 56807 299318 56835
rect 299346 56807 299380 56835
rect 299408 56807 299442 56835
rect 299470 56807 299518 56835
rect 299208 56773 299518 56807
rect 299208 56745 299256 56773
rect 299284 56745 299318 56773
rect 299346 56745 299380 56773
rect 299408 56745 299442 56773
rect 299470 56745 299518 56773
rect 299208 47959 299518 56745
rect 299208 47931 299256 47959
rect 299284 47931 299318 47959
rect 299346 47931 299380 47959
rect 299408 47931 299442 47959
rect 299470 47931 299518 47959
rect 299208 47897 299518 47931
rect 299208 47869 299256 47897
rect 299284 47869 299318 47897
rect 299346 47869 299380 47897
rect 299408 47869 299442 47897
rect 299470 47869 299518 47897
rect 299208 47835 299518 47869
rect 299208 47807 299256 47835
rect 299284 47807 299318 47835
rect 299346 47807 299380 47835
rect 299408 47807 299442 47835
rect 299470 47807 299518 47835
rect 299208 47773 299518 47807
rect 299208 47745 299256 47773
rect 299284 47745 299318 47773
rect 299346 47745 299380 47773
rect 299408 47745 299442 47773
rect 299470 47745 299518 47773
rect 299208 38959 299518 47745
rect 299208 38931 299256 38959
rect 299284 38931 299318 38959
rect 299346 38931 299380 38959
rect 299408 38931 299442 38959
rect 299470 38931 299518 38959
rect 299208 38897 299518 38931
rect 299208 38869 299256 38897
rect 299284 38869 299318 38897
rect 299346 38869 299380 38897
rect 299408 38869 299442 38897
rect 299470 38869 299518 38897
rect 299208 38835 299518 38869
rect 299208 38807 299256 38835
rect 299284 38807 299318 38835
rect 299346 38807 299380 38835
rect 299408 38807 299442 38835
rect 299470 38807 299518 38835
rect 299208 38773 299518 38807
rect 299208 38745 299256 38773
rect 299284 38745 299318 38773
rect 299346 38745 299380 38773
rect 299408 38745 299442 38773
rect 299470 38745 299518 38773
rect 299208 29959 299518 38745
rect 299208 29931 299256 29959
rect 299284 29931 299318 29959
rect 299346 29931 299380 29959
rect 299408 29931 299442 29959
rect 299470 29931 299518 29959
rect 299208 29897 299518 29931
rect 299208 29869 299256 29897
rect 299284 29869 299318 29897
rect 299346 29869 299380 29897
rect 299408 29869 299442 29897
rect 299470 29869 299518 29897
rect 299208 29835 299518 29869
rect 299208 29807 299256 29835
rect 299284 29807 299318 29835
rect 299346 29807 299380 29835
rect 299408 29807 299442 29835
rect 299470 29807 299518 29835
rect 299208 29773 299518 29807
rect 299208 29745 299256 29773
rect 299284 29745 299318 29773
rect 299346 29745 299380 29773
rect 299408 29745 299442 29773
rect 299470 29745 299518 29773
rect 299208 20959 299518 29745
rect 299208 20931 299256 20959
rect 299284 20931 299318 20959
rect 299346 20931 299380 20959
rect 299408 20931 299442 20959
rect 299470 20931 299518 20959
rect 299208 20897 299518 20931
rect 299208 20869 299256 20897
rect 299284 20869 299318 20897
rect 299346 20869 299380 20897
rect 299408 20869 299442 20897
rect 299470 20869 299518 20897
rect 299208 20835 299518 20869
rect 299208 20807 299256 20835
rect 299284 20807 299318 20835
rect 299346 20807 299380 20835
rect 299408 20807 299442 20835
rect 299470 20807 299518 20835
rect 299208 20773 299518 20807
rect 299208 20745 299256 20773
rect 299284 20745 299318 20773
rect 299346 20745 299380 20773
rect 299408 20745 299442 20773
rect 299470 20745 299518 20773
rect 299208 11959 299518 20745
rect 299208 11931 299256 11959
rect 299284 11931 299318 11959
rect 299346 11931 299380 11959
rect 299408 11931 299442 11959
rect 299470 11931 299518 11959
rect 299208 11897 299518 11931
rect 299208 11869 299256 11897
rect 299284 11869 299318 11897
rect 299346 11869 299380 11897
rect 299408 11869 299442 11897
rect 299470 11869 299518 11897
rect 299208 11835 299518 11869
rect 299208 11807 299256 11835
rect 299284 11807 299318 11835
rect 299346 11807 299380 11835
rect 299408 11807 299442 11835
rect 299470 11807 299518 11835
rect 299208 11773 299518 11807
rect 299208 11745 299256 11773
rect 299284 11745 299318 11773
rect 299346 11745 299380 11773
rect 299408 11745 299442 11773
rect 299470 11745 299518 11773
rect 299208 2959 299518 11745
rect 299208 2931 299256 2959
rect 299284 2931 299318 2959
rect 299346 2931 299380 2959
rect 299408 2931 299442 2959
rect 299470 2931 299518 2959
rect 299208 2897 299518 2931
rect 299208 2869 299256 2897
rect 299284 2869 299318 2897
rect 299346 2869 299380 2897
rect 299408 2869 299442 2897
rect 299470 2869 299518 2897
rect 299208 2835 299518 2869
rect 299208 2807 299256 2835
rect 299284 2807 299318 2835
rect 299346 2807 299380 2835
rect 299408 2807 299442 2835
rect 299470 2807 299518 2835
rect 299208 2773 299518 2807
rect 299208 2745 299256 2773
rect 299284 2745 299318 2773
rect 299346 2745 299380 2773
rect 299408 2745 299442 2773
rect 299470 2745 299518 2773
rect 299208 904 299518 2745
rect 299208 876 299256 904
rect 299284 876 299318 904
rect 299346 876 299380 904
rect 299408 876 299442 904
rect 299470 876 299518 904
rect 299208 842 299518 876
rect 299208 814 299256 842
rect 299284 814 299318 842
rect 299346 814 299380 842
rect 299408 814 299442 842
rect 299470 814 299518 842
rect 299208 780 299518 814
rect 299208 752 299256 780
rect 299284 752 299318 780
rect 299346 752 299380 780
rect 299408 752 299442 780
rect 299470 752 299518 780
rect 299208 718 299518 752
rect 299208 690 299256 718
rect 299284 690 299318 718
rect 299346 690 299380 718
rect 299408 690 299442 718
rect 299470 690 299518 718
rect 299208 642 299518 690
rect 299688 293959 299998 299456
rect 299688 293931 299736 293959
rect 299764 293931 299798 293959
rect 299826 293931 299860 293959
rect 299888 293931 299922 293959
rect 299950 293931 299998 293959
rect 299688 293897 299998 293931
rect 299688 293869 299736 293897
rect 299764 293869 299798 293897
rect 299826 293869 299860 293897
rect 299888 293869 299922 293897
rect 299950 293869 299998 293897
rect 299688 293835 299998 293869
rect 299688 293807 299736 293835
rect 299764 293807 299798 293835
rect 299826 293807 299860 293835
rect 299888 293807 299922 293835
rect 299950 293807 299998 293835
rect 299688 293773 299998 293807
rect 299688 293745 299736 293773
rect 299764 293745 299798 293773
rect 299826 293745 299860 293773
rect 299888 293745 299922 293773
rect 299950 293745 299998 293773
rect 299688 284959 299998 293745
rect 299688 284931 299736 284959
rect 299764 284931 299798 284959
rect 299826 284931 299860 284959
rect 299888 284931 299922 284959
rect 299950 284931 299998 284959
rect 299688 284897 299998 284931
rect 299688 284869 299736 284897
rect 299764 284869 299798 284897
rect 299826 284869 299860 284897
rect 299888 284869 299922 284897
rect 299950 284869 299998 284897
rect 299688 284835 299998 284869
rect 299688 284807 299736 284835
rect 299764 284807 299798 284835
rect 299826 284807 299860 284835
rect 299888 284807 299922 284835
rect 299950 284807 299998 284835
rect 299688 284773 299998 284807
rect 299688 284745 299736 284773
rect 299764 284745 299798 284773
rect 299826 284745 299860 284773
rect 299888 284745 299922 284773
rect 299950 284745 299998 284773
rect 299688 275959 299998 284745
rect 299688 275931 299736 275959
rect 299764 275931 299798 275959
rect 299826 275931 299860 275959
rect 299888 275931 299922 275959
rect 299950 275931 299998 275959
rect 299688 275897 299998 275931
rect 299688 275869 299736 275897
rect 299764 275869 299798 275897
rect 299826 275869 299860 275897
rect 299888 275869 299922 275897
rect 299950 275869 299998 275897
rect 299688 275835 299998 275869
rect 299688 275807 299736 275835
rect 299764 275807 299798 275835
rect 299826 275807 299860 275835
rect 299888 275807 299922 275835
rect 299950 275807 299998 275835
rect 299688 275773 299998 275807
rect 299688 275745 299736 275773
rect 299764 275745 299798 275773
rect 299826 275745 299860 275773
rect 299888 275745 299922 275773
rect 299950 275745 299998 275773
rect 299688 266959 299998 275745
rect 299688 266931 299736 266959
rect 299764 266931 299798 266959
rect 299826 266931 299860 266959
rect 299888 266931 299922 266959
rect 299950 266931 299998 266959
rect 299688 266897 299998 266931
rect 299688 266869 299736 266897
rect 299764 266869 299798 266897
rect 299826 266869 299860 266897
rect 299888 266869 299922 266897
rect 299950 266869 299998 266897
rect 299688 266835 299998 266869
rect 299688 266807 299736 266835
rect 299764 266807 299798 266835
rect 299826 266807 299860 266835
rect 299888 266807 299922 266835
rect 299950 266807 299998 266835
rect 299688 266773 299998 266807
rect 299688 266745 299736 266773
rect 299764 266745 299798 266773
rect 299826 266745 299860 266773
rect 299888 266745 299922 266773
rect 299950 266745 299998 266773
rect 299688 257959 299998 266745
rect 299688 257931 299736 257959
rect 299764 257931 299798 257959
rect 299826 257931 299860 257959
rect 299888 257931 299922 257959
rect 299950 257931 299998 257959
rect 299688 257897 299998 257931
rect 299688 257869 299736 257897
rect 299764 257869 299798 257897
rect 299826 257869 299860 257897
rect 299888 257869 299922 257897
rect 299950 257869 299998 257897
rect 299688 257835 299998 257869
rect 299688 257807 299736 257835
rect 299764 257807 299798 257835
rect 299826 257807 299860 257835
rect 299888 257807 299922 257835
rect 299950 257807 299998 257835
rect 299688 257773 299998 257807
rect 299688 257745 299736 257773
rect 299764 257745 299798 257773
rect 299826 257745 299860 257773
rect 299888 257745 299922 257773
rect 299950 257745 299998 257773
rect 299688 248959 299998 257745
rect 299688 248931 299736 248959
rect 299764 248931 299798 248959
rect 299826 248931 299860 248959
rect 299888 248931 299922 248959
rect 299950 248931 299998 248959
rect 299688 248897 299998 248931
rect 299688 248869 299736 248897
rect 299764 248869 299798 248897
rect 299826 248869 299860 248897
rect 299888 248869 299922 248897
rect 299950 248869 299998 248897
rect 299688 248835 299998 248869
rect 299688 248807 299736 248835
rect 299764 248807 299798 248835
rect 299826 248807 299860 248835
rect 299888 248807 299922 248835
rect 299950 248807 299998 248835
rect 299688 248773 299998 248807
rect 299688 248745 299736 248773
rect 299764 248745 299798 248773
rect 299826 248745 299860 248773
rect 299888 248745 299922 248773
rect 299950 248745 299998 248773
rect 299688 239959 299998 248745
rect 299688 239931 299736 239959
rect 299764 239931 299798 239959
rect 299826 239931 299860 239959
rect 299888 239931 299922 239959
rect 299950 239931 299998 239959
rect 299688 239897 299998 239931
rect 299688 239869 299736 239897
rect 299764 239869 299798 239897
rect 299826 239869 299860 239897
rect 299888 239869 299922 239897
rect 299950 239869 299998 239897
rect 299688 239835 299998 239869
rect 299688 239807 299736 239835
rect 299764 239807 299798 239835
rect 299826 239807 299860 239835
rect 299888 239807 299922 239835
rect 299950 239807 299998 239835
rect 299688 239773 299998 239807
rect 299688 239745 299736 239773
rect 299764 239745 299798 239773
rect 299826 239745 299860 239773
rect 299888 239745 299922 239773
rect 299950 239745 299998 239773
rect 299688 230959 299998 239745
rect 299688 230931 299736 230959
rect 299764 230931 299798 230959
rect 299826 230931 299860 230959
rect 299888 230931 299922 230959
rect 299950 230931 299998 230959
rect 299688 230897 299998 230931
rect 299688 230869 299736 230897
rect 299764 230869 299798 230897
rect 299826 230869 299860 230897
rect 299888 230869 299922 230897
rect 299950 230869 299998 230897
rect 299688 230835 299998 230869
rect 299688 230807 299736 230835
rect 299764 230807 299798 230835
rect 299826 230807 299860 230835
rect 299888 230807 299922 230835
rect 299950 230807 299998 230835
rect 299688 230773 299998 230807
rect 299688 230745 299736 230773
rect 299764 230745 299798 230773
rect 299826 230745 299860 230773
rect 299888 230745 299922 230773
rect 299950 230745 299998 230773
rect 299688 221959 299998 230745
rect 299688 221931 299736 221959
rect 299764 221931 299798 221959
rect 299826 221931 299860 221959
rect 299888 221931 299922 221959
rect 299950 221931 299998 221959
rect 299688 221897 299998 221931
rect 299688 221869 299736 221897
rect 299764 221869 299798 221897
rect 299826 221869 299860 221897
rect 299888 221869 299922 221897
rect 299950 221869 299998 221897
rect 299688 221835 299998 221869
rect 299688 221807 299736 221835
rect 299764 221807 299798 221835
rect 299826 221807 299860 221835
rect 299888 221807 299922 221835
rect 299950 221807 299998 221835
rect 299688 221773 299998 221807
rect 299688 221745 299736 221773
rect 299764 221745 299798 221773
rect 299826 221745 299860 221773
rect 299888 221745 299922 221773
rect 299950 221745 299998 221773
rect 299688 212959 299998 221745
rect 299688 212931 299736 212959
rect 299764 212931 299798 212959
rect 299826 212931 299860 212959
rect 299888 212931 299922 212959
rect 299950 212931 299998 212959
rect 299688 212897 299998 212931
rect 299688 212869 299736 212897
rect 299764 212869 299798 212897
rect 299826 212869 299860 212897
rect 299888 212869 299922 212897
rect 299950 212869 299998 212897
rect 299688 212835 299998 212869
rect 299688 212807 299736 212835
rect 299764 212807 299798 212835
rect 299826 212807 299860 212835
rect 299888 212807 299922 212835
rect 299950 212807 299998 212835
rect 299688 212773 299998 212807
rect 299688 212745 299736 212773
rect 299764 212745 299798 212773
rect 299826 212745 299860 212773
rect 299888 212745 299922 212773
rect 299950 212745 299998 212773
rect 299688 203959 299998 212745
rect 299688 203931 299736 203959
rect 299764 203931 299798 203959
rect 299826 203931 299860 203959
rect 299888 203931 299922 203959
rect 299950 203931 299998 203959
rect 299688 203897 299998 203931
rect 299688 203869 299736 203897
rect 299764 203869 299798 203897
rect 299826 203869 299860 203897
rect 299888 203869 299922 203897
rect 299950 203869 299998 203897
rect 299688 203835 299998 203869
rect 299688 203807 299736 203835
rect 299764 203807 299798 203835
rect 299826 203807 299860 203835
rect 299888 203807 299922 203835
rect 299950 203807 299998 203835
rect 299688 203773 299998 203807
rect 299688 203745 299736 203773
rect 299764 203745 299798 203773
rect 299826 203745 299860 203773
rect 299888 203745 299922 203773
rect 299950 203745 299998 203773
rect 299688 194959 299998 203745
rect 299688 194931 299736 194959
rect 299764 194931 299798 194959
rect 299826 194931 299860 194959
rect 299888 194931 299922 194959
rect 299950 194931 299998 194959
rect 299688 194897 299998 194931
rect 299688 194869 299736 194897
rect 299764 194869 299798 194897
rect 299826 194869 299860 194897
rect 299888 194869 299922 194897
rect 299950 194869 299998 194897
rect 299688 194835 299998 194869
rect 299688 194807 299736 194835
rect 299764 194807 299798 194835
rect 299826 194807 299860 194835
rect 299888 194807 299922 194835
rect 299950 194807 299998 194835
rect 299688 194773 299998 194807
rect 299688 194745 299736 194773
rect 299764 194745 299798 194773
rect 299826 194745 299860 194773
rect 299888 194745 299922 194773
rect 299950 194745 299998 194773
rect 299688 185959 299998 194745
rect 299688 185931 299736 185959
rect 299764 185931 299798 185959
rect 299826 185931 299860 185959
rect 299888 185931 299922 185959
rect 299950 185931 299998 185959
rect 299688 185897 299998 185931
rect 299688 185869 299736 185897
rect 299764 185869 299798 185897
rect 299826 185869 299860 185897
rect 299888 185869 299922 185897
rect 299950 185869 299998 185897
rect 299688 185835 299998 185869
rect 299688 185807 299736 185835
rect 299764 185807 299798 185835
rect 299826 185807 299860 185835
rect 299888 185807 299922 185835
rect 299950 185807 299998 185835
rect 299688 185773 299998 185807
rect 299688 185745 299736 185773
rect 299764 185745 299798 185773
rect 299826 185745 299860 185773
rect 299888 185745 299922 185773
rect 299950 185745 299998 185773
rect 299688 176959 299998 185745
rect 299688 176931 299736 176959
rect 299764 176931 299798 176959
rect 299826 176931 299860 176959
rect 299888 176931 299922 176959
rect 299950 176931 299998 176959
rect 299688 176897 299998 176931
rect 299688 176869 299736 176897
rect 299764 176869 299798 176897
rect 299826 176869 299860 176897
rect 299888 176869 299922 176897
rect 299950 176869 299998 176897
rect 299688 176835 299998 176869
rect 299688 176807 299736 176835
rect 299764 176807 299798 176835
rect 299826 176807 299860 176835
rect 299888 176807 299922 176835
rect 299950 176807 299998 176835
rect 299688 176773 299998 176807
rect 299688 176745 299736 176773
rect 299764 176745 299798 176773
rect 299826 176745 299860 176773
rect 299888 176745 299922 176773
rect 299950 176745 299998 176773
rect 299688 167959 299998 176745
rect 299688 167931 299736 167959
rect 299764 167931 299798 167959
rect 299826 167931 299860 167959
rect 299888 167931 299922 167959
rect 299950 167931 299998 167959
rect 299688 167897 299998 167931
rect 299688 167869 299736 167897
rect 299764 167869 299798 167897
rect 299826 167869 299860 167897
rect 299888 167869 299922 167897
rect 299950 167869 299998 167897
rect 299688 167835 299998 167869
rect 299688 167807 299736 167835
rect 299764 167807 299798 167835
rect 299826 167807 299860 167835
rect 299888 167807 299922 167835
rect 299950 167807 299998 167835
rect 299688 167773 299998 167807
rect 299688 167745 299736 167773
rect 299764 167745 299798 167773
rect 299826 167745 299860 167773
rect 299888 167745 299922 167773
rect 299950 167745 299998 167773
rect 299688 158959 299998 167745
rect 299688 158931 299736 158959
rect 299764 158931 299798 158959
rect 299826 158931 299860 158959
rect 299888 158931 299922 158959
rect 299950 158931 299998 158959
rect 299688 158897 299998 158931
rect 299688 158869 299736 158897
rect 299764 158869 299798 158897
rect 299826 158869 299860 158897
rect 299888 158869 299922 158897
rect 299950 158869 299998 158897
rect 299688 158835 299998 158869
rect 299688 158807 299736 158835
rect 299764 158807 299798 158835
rect 299826 158807 299860 158835
rect 299888 158807 299922 158835
rect 299950 158807 299998 158835
rect 299688 158773 299998 158807
rect 299688 158745 299736 158773
rect 299764 158745 299798 158773
rect 299826 158745 299860 158773
rect 299888 158745 299922 158773
rect 299950 158745 299998 158773
rect 299688 149959 299998 158745
rect 299688 149931 299736 149959
rect 299764 149931 299798 149959
rect 299826 149931 299860 149959
rect 299888 149931 299922 149959
rect 299950 149931 299998 149959
rect 299688 149897 299998 149931
rect 299688 149869 299736 149897
rect 299764 149869 299798 149897
rect 299826 149869 299860 149897
rect 299888 149869 299922 149897
rect 299950 149869 299998 149897
rect 299688 149835 299998 149869
rect 299688 149807 299736 149835
rect 299764 149807 299798 149835
rect 299826 149807 299860 149835
rect 299888 149807 299922 149835
rect 299950 149807 299998 149835
rect 299688 149773 299998 149807
rect 299688 149745 299736 149773
rect 299764 149745 299798 149773
rect 299826 149745 299860 149773
rect 299888 149745 299922 149773
rect 299950 149745 299998 149773
rect 299688 140959 299998 149745
rect 299688 140931 299736 140959
rect 299764 140931 299798 140959
rect 299826 140931 299860 140959
rect 299888 140931 299922 140959
rect 299950 140931 299998 140959
rect 299688 140897 299998 140931
rect 299688 140869 299736 140897
rect 299764 140869 299798 140897
rect 299826 140869 299860 140897
rect 299888 140869 299922 140897
rect 299950 140869 299998 140897
rect 299688 140835 299998 140869
rect 299688 140807 299736 140835
rect 299764 140807 299798 140835
rect 299826 140807 299860 140835
rect 299888 140807 299922 140835
rect 299950 140807 299998 140835
rect 299688 140773 299998 140807
rect 299688 140745 299736 140773
rect 299764 140745 299798 140773
rect 299826 140745 299860 140773
rect 299888 140745 299922 140773
rect 299950 140745 299998 140773
rect 299688 131959 299998 140745
rect 299688 131931 299736 131959
rect 299764 131931 299798 131959
rect 299826 131931 299860 131959
rect 299888 131931 299922 131959
rect 299950 131931 299998 131959
rect 299688 131897 299998 131931
rect 299688 131869 299736 131897
rect 299764 131869 299798 131897
rect 299826 131869 299860 131897
rect 299888 131869 299922 131897
rect 299950 131869 299998 131897
rect 299688 131835 299998 131869
rect 299688 131807 299736 131835
rect 299764 131807 299798 131835
rect 299826 131807 299860 131835
rect 299888 131807 299922 131835
rect 299950 131807 299998 131835
rect 299688 131773 299998 131807
rect 299688 131745 299736 131773
rect 299764 131745 299798 131773
rect 299826 131745 299860 131773
rect 299888 131745 299922 131773
rect 299950 131745 299998 131773
rect 299688 122959 299998 131745
rect 299688 122931 299736 122959
rect 299764 122931 299798 122959
rect 299826 122931 299860 122959
rect 299888 122931 299922 122959
rect 299950 122931 299998 122959
rect 299688 122897 299998 122931
rect 299688 122869 299736 122897
rect 299764 122869 299798 122897
rect 299826 122869 299860 122897
rect 299888 122869 299922 122897
rect 299950 122869 299998 122897
rect 299688 122835 299998 122869
rect 299688 122807 299736 122835
rect 299764 122807 299798 122835
rect 299826 122807 299860 122835
rect 299888 122807 299922 122835
rect 299950 122807 299998 122835
rect 299688 122773 299998 122807
rect 299688 122745 299736 122773
rect 299764 122745 299798 122773
rect 299826 122745 299860 122773
rect 299888 122745 299922 122773
rect 299950 122745 299998 122773
rect 299688 113959 299998 122745
rect 299688 113931 299736 113959
rect 299764 113931 299798 113959
rect 299826 113931 299860 113959
rect 299888 113931 299922 113959
rect 299950 113931 299998 113959
rect 299688 113897 299998 113931
rect 299688 113869 299736 113897
rect 299764 113869 299798 113897
rect 299826 113869 299860 113897
rect 299888 113869 299922 113897
rect 299950 113869 299998 113897
rect 299688 113835 299998 113869
rect 299688 113807 299736 113835
rect 299764 113807 299798 113835
rect 299826 113807 299860 113835
rect 299888 113807 299922 113835
rect 299950 113807 299998 113835
rect 299688 113773 299998 113807
rect 299688 113745 299736 113773
rect 299764 113745 299798 113773
rect 299826 113745 299860 113773
rect 299888 113745 299922 113773
rect 299950 113745 299998 113773
rect 299688 104959 299998 113745
rect 299688 104931 299736 104959
rect 299764 104931 299798 104959
rect 299826 104931 299860 104959
rect 299888 104931 299922 104959
rect 299950 104931 299998 104959
rect 299688 104897 299998 104931
rect 299688 104869 299736 104897
rect 299764 104869 299798 104897
rect 299826 104869 299860 104897
rect 299888 104869 299922 104897
rect 299950 104869 299998 104897
rect 299688 104835 299998 104869
rect 299688 104807 299736 104835
rect 299764 104807 299798 104835
rect 299826 104807 299860 104835
rect 299888 104807 299922 104835
rect 299950 104807 299998 104835
rect 299688 104773 299998 104807
rect 299688 104745 299736 104773
rect 299764 104745 299798 104773
rect 299826 104745 299860 104773
rect 299888 104745 299922 104773
rect 299950 104745 299998 104773
rect 299688 95959 299998 104745
rect 299688 95931 299736 95959
rect 299764 95931 299798 95959
rect 299826 95931 299860 95959
rect 299888 95931 299922 95959
rect 299950 95931 299998 95959
rect 299688 95897 299998 95931
rect 299688 95869 299736 95897
rect 299764 95869 299798 95897
rect 299826 95869 299860 95897
rect 299888 95869 299922 95897
rect 299950 95869 299998 95897
rect 299688 95835 299998 95869
rect 299688 95807 299736 95835
rect 299764 95807 299798 95835
rect 299826 95807 299860 95835
rect 299888 95807 299922 95835
rect 299950 95807 299998 95835
rect 299688 95773 299998 95807
rect 299688 95745 299736 95773
rect 299764 95745 299798 95773
rect 299826 95745 299860 95773
rect 299888 95745 299922 95773
rect 299950 95745 299998 95773
rect 299688 86959 299998 95745
rect 299688 86931 299736 86959
rect 299764 86931 299798 86959
rect 299826 86931 299860 86959
rect 299888 86931 299922 86959
rect 299950 86931 299998 86959
rect 299688 86897 299998 86931
rect 299688 86869 299736 86897
rect 299764 86869 299798 86897
rect 299826 86869 299860 86897
rect 299888 86869 299922 86897
rect 299950 86869 299998 86897
rect 299688 86835 299998 86869
rect 299688 86807 299736 86835
rect 299764 86807 299798 86835
rect 299826 86807 299860 86835
rect 299888 86807 299922 86835
rect 299950 86807 299998 86835
rect 299688 86773 299998 86807
rect 299688 86745 299736 86773
rect 299764 86745 299798 86773
rect 299826 86745 299860 86773
rect 299888 86745 299922 86773
rect 299950 86745 299998 86773
rect 299688 77959 299998 86745
rect 299688 77931 299736 77959
rect 299764 77931 299798 77959
rect 299826 77931 299860 77959
rect 299888 77931 299922 77959
rect 299950 77931 299998 77959
rect 299688 77897 299998 77931
rect 299688 77869 299736 77897
rect 299764 77869 299798 77897
rect 299826 77869 299860 77897
rect 299888 77869 299922 77897
rect 299950 77869 299998 77897
rect 299688 77835 299998 77869
rect 299688 77807 299736 77835
rect 299764 77807 299798 77835
rect 299826 77807 299860 77835
rect 299888 77807 299922 77835
rect 299950 77807 299998 77835
rect 299688 77773 299998 77807
rect 299688 77745 299736 77773
rect 299764 77745 299798 77773
rect 299826 77745 299860 77773
rect 299888 77745 299922 77773
rect 299950 77745 299998 77773
rect 299688 68959 299998 77745
rect 299688 68931 299736 68959
rect 299764 68931 299798 68959
rect 299826 68931 299860 68959
rect 299888 68931 299922 68959
rect 299950 68931 299998 68959
rect 299688 68897 299998 68931
rect 299688 68869 299736 68897
rect 299764 68869 299798 68897
rect 299826 68869 299860 68897
rect 299888 68869 299922 68897
rect 299950 68869 299998 68897
rect 299688 68835 299998 68869
rect 299688 68807 299736 68835
rect 299764 68807 299798 68835
rect 299826 68807 299860 68835
rect 299888 68807 299922 68835
rect 299950 68807 299998 68835
rect 299688 68773 299998 68807
rect 299688 68745 299736 68773
rect 299764 68745 299798 68773
rect 299826 68745 299860 68773
rect 299888 68745 299922 68773
rect 299950 68745 299998 68773
rect 299688 59959 299998 68745
rect 299688 59931 299736 59959
rect 299764 59931 299798 59959
rect 299826 59931 299860 59959
rect 299888 59931 299922 59959
rect 299950 59931 299998 59959
rect 299688 59897 299998 59931
rect 299688 59869 299736 59897
rect 299764 59869 299798 59897
rect 299826 59869 299860 59897
rect 299888 59869 299922 59897
rect 299950 59869 299998 59897
rect 299688 59835 299998 59869
rect 299688 59807 299736 59835
rect 299764 59807 299798 59835
rect 299826 59807 299860 59835
rect 299888 59807 299922 59835
rect 299950 59807 299998 59835
rect 299688 59773 299998 59807
rect 299688 59745 299736 59773
rect 299764 59745 299798 59773
rect 299826 59745 299860 59773
rect 299888 59745 299922 59773
rect 299950 59745 299998 59773
rect 299688 50959 299998 59745
rect 299688 50931 299736 50959
rect 299764 50931 299798 50959
rect 299826 50931 299860 50959
rect 299888 50931 299922 50959
rect 299950 50931 299998 50959
rect 299688 50897 299998 50931
rect 299688 50869 299736 50897
rect 299764 50869 299798 50897
rect 299826 50869 299860 50897
rect 299888 50869 299922 50897
rect 299950 50869 299998 50897
rect 299688 50835 299998 50869
rect 299688 50807 299736 50835
rect 299764 50807 299798 50835
rect 299826 50807 299860 50835
rect 299888 50807 299922 50835
rect 299950 50807 299998 50835
rect 299688 50773 299998 50807
rect 299688 50745 299736 50773
rect 299764 50745 299798 50773
rect 299826 50745 299860 50773
rect 299888 50745 299922 50773
rect 299950 50745 299998 50773
rect 299688 41959 299998 50745
rect 299688 41931 299736 41959
rect 299764 41931 299798 41959
rect 299826 41931 299860 41959
rect 299888 41931 299922 41959
rect 299950 41931 299998 41959
rect 299688 41897 299998 41931
rect 299688 41869 299736 41897
rect 299764 41869 299798 41897
rect 299826 41869 299860 41897
rect 299888 41869 299922 41897
rect 299950 41869 299998 41897
rect 299688 41835 299998 41869
rect 299688 41807 299736 41835
rect 299764 41807 299798 41835
rect 299826 41807 299860 41835
rect 299888 41807 299922 41835
rect 299950 41807 299998 41835
rect 299688 41773 299998 41807
rect 299688 41745 299736 41773
rect 299764 41745 299798 41773
rect 299826 41745 299860 41773
rect 299888 41745 299922 41773
rect 299950 41745 299998 41773
rect 299688 32959 299998 41745
rect 299688 32931 299736 32959
rect 299764 32931 299798 32959
rect 299826 32931 299860 32959
rect 299888 32931 299922 32959
rect 299950 32931 299998 32959
rect 299688 32897 299998 32931
rect 299688 32869 299736 32897
rect 299764 32869 299798 32897
rect 299826 32869 299860 32897
rect 299888 32869 299922 32897
rect 299950 32869 299998 32897
rect 299688 32835 299998 32869
rect 299688 32807 299736 32835
rect 299764 32807 299798 32835
rect 299826 32807 299860 32835
rect 299888 32807 299922 32835
rect 299950 32807 299998 32835
rect 299688 32773 299998 32807
rect 299688 32745 299736 32773
rect 299764 32745 299798 32773
rect 299826 32745 299860 32773
rect 299888 32745 299922 32773
rect 299950 32745 299998 32773
rect 299688 23959 299998 32745
rect 299688 23931 299736 23959
rect 299764 23931 299798 23959
rect 299826 23931 299860 23959
rect 299888 23931 299922 23959
rect 299950 23931 299998 23959
rect 299688 23897 299998 23931
rect 299688 23869 299736 23897
rect 299764 23869 299798 23897
rect 299826 23869 299860 23897
rect 299888 23869 299922 23897
rect 299950 23869 299998 23897
rect 299688 23835 299998 23869
rect 299688 23807 299736 23835
rect 299764 23807 299798 23835
rect 299826 23807 299860 23835
rect 299888 23807 299922 23835
rect 299950 23807 299998 23835
rect 299688 23773 299998 23807
rect 299688 23745 299736 23773
rect 299764 23745 299798 23773
rect 299826 23745 299860 23773
rect 299888 23745 299922 23773
rect 299950 23745 299998 23773
rect 299688 14959 299998 23745
rect 299688 14931 299736 14959
rect 299764 14931 299798 14959
rect 299826 14931 299860 14959
rect 299888 14931 299922 14959
rect 299950 14931 299998 14959
rect 299688 14897 299998 14931
rect 299688 14869 299736 14897
rect 299764 14869 299798 14897
rect 299826 14869 299860 14897
rect 299888 14869 299922 14897
rect 299950 14869 299998 14897
rect 299688 14835 299998 14869
rect 299688 14807 299736 14835
rect 299764 14807 299798 14835
rect 299826 14807 299860 14835
rect 299888 14807 299922 14835
rect 299950 14807 299998 14835
rect 299688 14773 299998 14807
rect 299688 14745 299736 14773
rect 299764 14745 299798 14773
rect 299826 14745 299860 14773
rect 299888 14745 299922 14773
rect 299950 14745 299998 14773
rect 299688 5959 299998 14745
rect 299688 5931 299736 5959
rect 299764 5931 299798 5959
rect 299826 5931 299860 5959
rect 299888 5931 299922 5959
rect 299950 5931 299998 5959
rect 299688 5897 299998 5931
rect 299688 5869 299736 5897
rect 299764 5869 299798 5897
rect 299826 5869 299860 5897
rect 299888 5869 299922 5897
rect 299950 5869 299998 5897
rect 299688 5835 299998 5869
rect 299688 5807 299736 5835
rect 299764 5807 299798 5835
rect 299826 5807 299860 5835
rect 299888 5807 299922 5835
rect 299950 5807 299998 5835
rect 299688 5773 299998 5807
rect 299688 5745 299736 5773
rect 299764 5745 299798 5773
rect 299826 5745 299860 5773
rect 299888 5745 299922 5773
rect 299950 5745 299998 5773
rect 292389 396 292437 424
rect 292465 396 292499 424
rect 292527 396 292561 424
rect 292589 396 292623 424
rect 292651 396 292699 424
rect 292389 362 292699 396
rect 292389 334 292437 362
rect 292465 334 292499 362
rect 292527 334 292561 362
rect 292589 334 292623 362
rect 292651 334 292699 362
rect 292389 300 292699 334
rect 292389 272 292437 300
rect 292465 272 292499 300
rect 292527 272 292561 300
rect 292589 272 292623 300
rect 292651 272 292699 300
rect 292389 238 292699 272
rect 292389 210 292437 238
rect 292465 210 292499 238
rect 292527 210 292561 238
rect 292589 210 292623 238
rect 292651 210 292699 238
rect 292389 162 292699 210
rect 299688 424 299998 5745
rect 299688 396 299736 424
rect 299764 396 299798 424
rect 299826 396 299860 424
rect 299888 396 299922 424
rect 299950 396 299998 424
rect 299688 362 299998 396
rect 299688 334 299736 362
rect 299764 334 299798 362
rect 299826 334 299860 362
rect 299888 334 299922 362
rect 299950 334 299998 362
rect 299688 300 299998 334
rect 299688 272 299736 300
rect 299764 272 299798 300
rect 299826 272 299860 300
rect 299888 272 299922 300
rect 299950 272 299998 300
rect 299688 238 299998 272
rect 299688 210 299736 238
rect 299764 210 299798 238
rect 299826 210 299860 238
rect 299888 210 299922 238
rect 299950 210 299998 238
rect 299688 162 299998 210
<< via4 >>
rect 42 299642 70 299670
rect 104 299642 132 299670
rect 166 299642 194 299670
rect 228 299642 256 299670
rect 42 299580 70 299608
rect 104 299580 132 299608
rect 166 299580 194 299608
rect 228 299580 256 299608
rect 42 299518 70 299546
rect 104 299518 132 299546
rect 166 299518 194 299546
rect 228 299518 256 299546
rect 42 299456 70 299484
rect 104 299456 132 299484
rect 166 299456 194 299484
rect 228 299456 256 299484
rect 42 293931 70 293959
rect 104 293931 132 293959
rect 166 293931 194 293959
rect 228 293931 256 293959
rect 42 293869 70 293897
rect 104 293869 132 293897
rect 166 293869 194 293897
rect 228 293869 256 293897
rect 42 293807 70 293835
rect 104 293807 132 293835
rect 166 293807 194 293835
rect 228 293807 256 293835
rect 42 293745 70 293773
rect 104 293745 132 293773
rect 166 293745 194 293773
rect 228 293745 256 293773
rect 42 284931 70 284959
rect 104 284931 132 284959
rect 166 284931 194 284959
rect 228 284931 256 284959
rect 42 284869 70 284897
rect 104 284869 132 284897
rect 166 284869 194 284897
rect 228 284869 256 284897
rect 42 284807 70 284835
rect 104 284807 132 284835
rect 166 284807 194 284835
rect 228 284807 256 284835
rect 42 284745 70 284773
rect 104 284745 132 284773
rect 166 284745 194 284773
rect 228 284745 256 284773
rect 42 275931 70 275959
rect 104 275931 132 275959
rect 166 275931 194 275959
rect 228 275931 256 275959
rect 42 275869 70 275897
rect 104 275869 132 275897
rect 166 275869 194 275897
rect 228 275869 256 275897
rect 42 275807 70 275835
rect 104 275807 132 275835
rect 166 275807 194 275835
rect 228 275807 256 275835
rect 42 275745 70 275773
rect 104 275745 132 275773
rect 166 275745 194 275773
rect 228 275745 256 275773
rect 42 266931 70 266959
rect 104 266931 132 266959
rect 166 266931 194 266959
rect 228 266931 256 266959
rect 42 266869 70 266897
rect 104 266869 132 266897
rect 166 266869 194 266897
rect 228 266869 256 266897
rect 42 266807 70 266835
rect 104 266807 132 266835
rect 166 266807 194 266835
rect 228 266807 256 266835
rect 42 266745 70 266773
rect 104 266745 132 266773
rect 166 266745 194 266773
rect 228 266745 256 266773
rect 42 257931 70 257959
rect 104 257931 132 257959
rect 166 257931 194 257959
rect 228 257931 256 257959
rect 42 257869 70 257897
rect 104 257869 132 257897
rect 166 257869 194 257897
rect 228 257869 256 257897
rect 42 257807 70 257835
rect 104 257807 132 257835
rect 166 257807 194 257835
rect 228 257807 256 257835
rect 42 257745 70 257773
rect 104 257745 132 257773
rect 166 257745 194 257773
rect 228 257745 256 257773
rect 42 248931 70 248959
rect 104 248931 132 248959
rect 166 248931 194 248959
rect 228 248931 256 248959
rect 42 248869 70 248897
rect 104 248869 132 248897
rect 166 248869 194 248897
rect 228 248869 256 248897
rect 42 248807 70 248835
rect 104 248807 132 248835
rect 166 248807 194 248835
rect 228 248807 256 248835
rect 42 248745 70 248773
rect 104 248745 132 248773
rect 166 248745 194 248773
rect 228 248745 256 248773
rect 42 239931 70 239959
rect 104 239931 132 239959
rect 166 239931 194 239959
rect 228 239931 256 239959
rect 42 239869 70 239897
rect 104 239869 132 239897
rect 166 239869 194 239897
rect 228 239869 256 239897
rect 42 239807 70 239835
rect 104 239807 132 239835
rect 166 239807 194 239835
rect 228 239807 256 239835
rect 42 239745 70 239773
rect 104 239745 132 239773
rect 166 239745 194 239773
rect 228 239745 256 239773
rect 42 230931 70 230959
rect 104 230931 132 230959
rect 166 230931 194 230959
rect 228 230931 256 230959
rect 42 230869 70 230897
rect 104 230869 132 230897
rect 166 230869 194 230897
rect 228 230869 256 230897
rect 42 230807 70 230835
rect 104 230807 132 230835
rect 166 230807 194 230835
rect 228 230807 256 230835
rect 42 230745 70 230773
rect 104 230745 132 230773
rect 166 230745 194 230773
rect 228 230745 256 230773
rect 42 221931 70 221959
rect 104 221931 132 221959
rect 166 221931 194 221959
rect 228 221931 256 221959
rect 42 221869 70 221897
rect 104 221869 132 221897
rect 166 221869 194 221897
rect 228 221869 256 221897
rect 42 221807 70 221835
rect 104 221807 132 221835
rect 166 221807 194 221835
rect 228 221807 256 221835
rect 42 221745 70 221773
rect 104 221745 132 221773
rect 166 221745 194 221773
rect 228 221745 256 221773
rect 42 212931 70 212959
rect 104 212931 132 212959
rect 166 212931 194 212959
rect 228 212931 256 212959
rect 42 212869 70 212897
rect 104 212869 132 212897
rect 166 212869 194 212897
rect 228 212869 256 212897
rect 42 212807 70 212835
rect 104 212807 132 212835
rect 166 212807 194 212835
rect 228 212807 256 212835
rect 42 212745 70 212773
rect 104 212745 132 212773
rect 166 212745 194 212773
rect 228 212745 256 212773
rect 42 203931 70 203959
rect 104 203931 132 203959
rect 166 203931 194 203959
rect 228 203931 256 203959
rect 42 203869 70 203897
rect 104 203869 132 203897
rect 166 203869 194 203897
rect 228 203869 256 203897
rect 42 203807 70 203835
rect 104 203807 132 203835
rect 166 203807 194 203835
rect 228 203807 256 203835
rect 42 203745 70 203773
rect 104 203745 132 203773
rect 166 203745 194 203773
rect 228 203745 256 203773
rect 42 194931 70 194959
rect 104 194931 132 194959
rect 166 194931 194 194959
rect 228 194931 256 194959
rect 42 194869 70 194897
rect 104 194869 132 194897
rect 166 194869 194 194897
rect 228 194869 256 194897
rect 42 194807 70 194835
rect 104 194807 132 194835
rect 166 194807 194 194835
rect 228 194807 256 194835
rect 42 194745 70 194773
rect 104 194745 132 194773
rect 166 194745 194 194773
rect 228 194745 256 194773
rect 42 185931 70 185959
rect 104 185931 132 185959
rect 166 185931 194 185959
rect 228 185931 256 185959
rect 42 185869 70 185897
rect 104 185869 132 185897
rect 166 185869 194 185897
rect 228 185869 256 185897
rect 42 185807 70 185835
rect 104 185807 132 185835
rect 166 185807 194 185835
rect 228 185807 256 185835
rect 42 185745 70 185773
rect 104 185745 132 185773
rect 166 185745 194 185773
rect 228 185745 256 185773
rect 42 176931 70 176959
rect 104 176931 132 176959
rect 166 176931 194 176959
rect 228 176931 256 176959
rect 42 176869 70 176897
rect 104 176869 132 176897
rect 166 176869 194 176897
rect 228 176869 256 176897
rect 42 176807 70 176835
rect 104 176807 132 176835
rect 166 176807 194 176835
rect 228 176807 256 176835
rect 42 176745 70 176773
rect 104 176745 132 176773
rect 166 176745 194 176773
rect 228 176745 256 176773
rect 42 167931 70 167959
rect 104 167931 132 167959
rect 166 167931 194 167959
rect 228 167931 256 167959
rect 42 167869 70 167897
rect 104 167869 132 167897
rect 166 167869 194 167897
rect 228 167869 256 167897
rect 42 167807 70 167835
rect 104 167807 132 167835
rect 166 167807 194 167835
rect 228 167807 256 167835
rect 42 167745 70 167773
rect 104 167745 132 167773
rect 166 167745 194 167773
rect 228 167745 256 167773
rect 42 158931 70 158959
rect 104 158931 132 158959
rect 166 158931 194 158959
rect 228 158931 256 158959
rect 42 158869 70 158897
rect 104 158869 132 158897
rect 166 158869 194 158897
rect 228 158869 256 158897
rect 42 158807 70 158835
rect 104 158807 132 158835
rect 166 158807 194 158835
rect 228 158807 256 158835
rect 42 158745 70 158773
rect 104 158745 132 158773
rect 166 158745 194 158773
rect 228 158745 256 158773
rect 42 149931 70 149959
rect 104 149931 132 149959
rect 166 149931 194 149959
rect 228 149931 256 149959
rect 42 149869 70 149897
rect 104 149869 132 149897
rect 166 149869 194 149897
rect 228 149869 256 149897
rect 42 149807 70 149835
rect 104 149807 132 149835
rect 166 149807 194 149835
rect 228 149807 256 149835
rect 42 149745 70 149773
rect 104 149745 132 149773
rect 166 149745 194 149773
rect 228 149745 256 149773
rect 42 140931 70 140959
rect 104 140931 132 140959
rect 166 140931 194 140959
rect 228 140931 256 140959
rect 42 140869 70 140897
rect 104 140869 132 140897
rect 166 140869 194 140897
rect 228 140869 256 140897
rect 42 140807 70 140835
rect 104 140807 132 140835
rect 166 140807 194 140835
rect 228 140807 256 140835
rect 42 140745 70 140773
rect 104 140745 132 140773
rect 166 140745 194 140773
rect 228 140745 256 140773
rect 42 131931 70 131959
rect 104 131931 132 131959
rect 166 131931 194 131959
rect 228 131931 256 131959
rect 42 131869 70 131897
rect 104 131869 132 131897
rect 166 131869 194 131897
rect 228 131869 256 131897
rect 42 131807 70 131835
rect 104 131807 132 131835
rect 166 131807 194 131835
rect 228 131807 256 131835
rect 42 131745 70 131773
rect 104 131745 132 131773
rect 166 131745 194 131773
rect 228 131745 256 131773
rect 42 122931 70 122959
rect 104 122931 132 122959
rect 166 122931 194 122959
rect 228 122931 256 122959
rect 42 122869 70 122897
rect 104 122869 132 122897
rect 166 122869 194 122897
rect 228 122869 256 122897
rect 42 122807 70 122835
rect 104 122807 132 122835
rect 166 122807 194 122835
rect 228 122807 256 122835
rect 42 122745 70 122773
rect 104 122745 132 122773
rect 166 122745 194 122773
rect 228 122745 256 122773
rect 42 113931 70 113959
rect 104 113931 132 113959
rect 166 113931 194 113959
rect 228 113931 256 113959
rect 42 113869 70 113897
rect 104 113869 132 113897
rect 166 113869 194 113897
rect 228 113869 256 113897
rect 42 113807 70 113835
rect 104 113807 132 113835
rect 166 113807 194 113835
rect 228 113807 256 113835
rect 42 113745 70 113773
rect 104 113745 132 113773
rect 166 113745 194 113773
rect 228 113745 256 113773
rect 42 104931 70 104959
rect 104 104931 132 104959
rect 166 104931 194 104959
rect 228 104931 256 104959
rect 42 104869 70 104897
rect 104 104869 132 104897
rect 166 104869 194 104897
rect 228 104869 256 104897
rect 42 104807 70 104835
rect 104 104807 132 104835
rect 166 104807 194 104835
rect 228 104807 256 104835
rect 42 104745 70 104773
rect 104 104745 132 104773
rect 166 104745 194 104773
rect 228 104745 256 104773
rect 42 95931 70 95959
rect 104 95931 132 95959
rect 166 95931 194 95959
rect 228 95931 256 95959
rect 42 95869 70 95897
rect 104 95869 132 95897
rect 166 95869 194 95897
rect 228 95869 256 95897
rect 42 95807 70 95835
rect 104 95807 132 95835
rect 166 95807 194 95835
rect 228 95807 256 95835
rect 42 95745 70 95773
rect 104 95745 132 95773
rect 166 95745 194 95773
rect 228 95745 256 95773
rect 42 86931 70 86959
rect 104 86931 132 86959
rect 166 86931 194 86959
rect 228 86931 256 86959
rect 42 86869 70 86897
rect 104 86869 132 86897
rect 166 86869 194 86897
rect 228 86869 256 86897
rect 42 86807 70 86835
rect 104 86807 132 86835
rect 166 86807 194 86835
rect 228 86807 256 86835
rect 42 86745 70 86773
rect 104 86745 132 86773
rect 166 86745 194 86773
rect 228 86745 256 86773
rect 42 77931 70 77959
rect 104 77931 132 77959
rect 166 77931 194 77959
rect 228 77931 256 77959
rect 42 77869 70 77897
rect 104 77869 132 77897
rect 166 77869 194 77897
rect 228 77869 256 77897
rect 42 77807 70 77835
rect 104 77807 132 77835
rect 166 77807 194 77835
rect 228 77807 256 77835
rect 42 77745 70 77773
rect 104 77745 132 77773
rect 166 77745 194 77773
rect 228 77745 256 77773
rect 42 68931 70 68959
rect 104 68931 132 68959
rect 166 68931 194 68959
rect 228 68931 256 68959
rect 42 68869 70 68897
rect 104 68869 132 68897
rect 166 68869 194 68897
rect 228 68869 256 68897
rect 42 68807 70 68835
rect 104 68807 132 68835
rect 166 68807 194 68835
rect 228 68807 256 68835
rect 42 68745 70 68773
rect 104 68745 132 68773
rect 166 68745 194 68773
rect 228 68745 256 68773
rect 42 59931 70 59959
rect 104 59931 132 59959
rect 166 59931 194 59959
rect 228 59931 256 59959
rect 42 59869 70 59897
rect 104 59869 132 59897
rect 166 59869 194 59897
rect 228 59869 256 59897
rect 42 59807 70 59835
rect 104 59807 132 59835
rect 166 59807 194 59835
rect 228 59807 256 59835
rect 42 59745 70 59773
rect 104 59745 132 59773
rect 166 59745 194 59773
rect 228 59745 256 59773
rect 42 50931 70 50959
rect 104 50931 132 50959
rect 166 50931 194 50959
rect 228 50931 256 50959
rect 42 50869 70 50897
rect 104 50869 132 50897
rect 166 50869 194 50897
rect 228 50869 256 50897
rect 42 50807 70 50835
rect 104 50807 132 50835
rect 166 50807 194 50835
rect 228 50807 256 50835
rect 42 50745 70 50773
rect 104 50745 132 50773
rect 166 50745 194 50773
rect 228 50745 256 50773
rect 42 41931 70 41959
rect 104 41931 132 41959
rect 166 41931 194 41959
rect 228 41931 256 41959
rect 42 41869 70 41897
rect 104 41869 132 41897
rect 166 41869 194 41897
rect 228 41869 256 41897
rect 42 41807 70 41835
rect 104 41807 132 41835
rect 166 41807 194 41835
rect 228 41807 256 41835
rect 42 41745 70 41773
rect 104 41745 132 41773
rect 166 41745 194 41773
rect 228 41745 256 41773
rect 42 32931 70 32959
rect 104 32931 132 32959
rect 166 32931 194 32959
rect 228 32931 256 32959
rect 42 32869 70 32897
rect 104 32869 132 32897
rect 166 32869 194 32897
rect 228 32869 256 32897
rect 42 32807 70 32835
rect 104 32807 132 32835
rect 166 32807 194 32835
rect 228 32807 256 32835
rect 42 32745 70 32773
rect 104 32745 132 32773
rect 166 32745 194 32773
rect 228 32745 256 32773
rect 42 23931 70 23959
rect 104 23931 132 23959
rect 166 23931 194 23959
rect 228 23931 256 23959
rect 42 23869 70 23897
rect 104 23869 132 23897
rect 166 23869 194 23897
rect 228 23869 256 23897
rect 42 23807 70 23835
rect 104 23807 132 23835
rect 166 23807 194 23835
rect 228 23807 256 23835
rect 42 23745 70 23773
rect 104 23745 132 23773
rect 166 23745 194 23773
rect 228 23745 256 23773
rect 42 14931 70 14959
rect 104 14931 132 14959
rect 166 14931 194 14959
rect 228 14931 256 14959
rect 42 14869 70 14897
rect 104 14869 132 14897
rect 166 14869 194 14897
rect 228 14869 256 14897
rect 42 14807 70 14835
rect 104 14807 132 14835
rect 166 14807 194 14835
rect 228 14807 256 14835
rect 42 14745 70 14773
rect 104 14745 132 14773
rect 166 14745 194 14773
rect 228 14745 256 14773
rect 42 5931 70 5959
rect 104 5931 132 5959
rect 166 5931 194 5959
rect 228 5931 256 5959
rect 42 5869 70 5897
rect 104 5869 132 5897
rect 166 5869 194 5897
rect 228 5869 256 5897
rect 42 5807 70 5835
rect 104 5807 132 5835
rect 166 5807 194 5835
rect 228 5807 256 5835
rect 42 5745 70 5773
rect 104 5745 132 5773
rect 166 5745 194 5773
rect 228 5745 256 5773
rect 522 299162 550 299190
rect 584 299162 612 299190
rect 646 299162 674 299190
rect 708 299162 736 299190
rect 522 299100 550 299128
rect 584 299100 612 299128
rect 646 299100 674 299128
rect 708 299100 736 299128
rect 522 299038 550 299066
rect 584 299038 612 299066
rect 646 299038 674 299066
rect 708 299038 736 299066
rect 522 298976 550 299004
rect 584 298976 612 299004
rect 646 298976 674 299004
rect 708 298976 736 299004
rect 522 290931 550 290959
rect 584 290931 612 290959
rect 646 290931 674 290959
rect 708 290931 736 290959
rect 522 290869 550 290897
rect 584 290869 612 290897
rect 646 290869 674 290897
rect 708 290869 736 290897
rect 522 290807 550 290835
rect 584 290807 612 290835
rect 646 290807 674 290835
rect 708 290807 736 290835
rect 522 290745 550 290773
rect 584 290745 612 290773
rect 646 290745 674 290773
rect 708 290745 736 290773
rect 522 281931 550 281959
rect 584 281931 612 281959
rect 646 281931 674 281959
rect 708 281931 736 281959
rect 522 281869 550 281897
rect 584 281869 612 281897
rect 646 281869 674 281897
rect 708 281869 736 281897
rect 522 281807 550 281835
rect 584 281807 612 281835
rect 646 281807 674 281835
rect 708 281807 736 281835
rect 522 281745 550 281773
rect 584 281745 612 281773
rect 646 281745 674 281773
rect 708 281745 736 281773
rect 522 272931 550 272959
rect 584 272931 612 272959
rect 646 272931 674 272959
rect 708 272931 736 272959
rect 522 272869 550 272897
rect 584 272869 612 272897
rect 646 272869 674 272897
rect 708 272869 736 272897
rect 522 272807 550 272835
rect 584 272807 612 272835
rect 646 272807 674 272835
rect 708 272807 736 272835
rect 522 272745 550 272773
rect 584 272745 612 272773
rect 646 272745 674 272773
rect 708 272745 736 272773
rect 522 263931 550 263959
rect 584 263931 612 263959
rect 646 263931 674 263959
rect 708 263931 736 263959
rect 522 263869 550 263897
rect 584 263869 612 263897
rect 646 263869 674 263897
rect 708 263869 736 263897
rect 522 263807 550 263835
rect 584 263807 612 263835
rect 646 263807 674 263835
rect 708 263807 736 263835
rect 522 263745 550 263773
rect 584 263745 612 263773
rect 646 263745 674 263773
rect 708 263745 736 263773
rect 522 254931 550 254959
rect 584 254931 612 254959
rect 646 254931 674 254959
rect 708 254931 736 254959
rect 522 254869 550 254897
rect 584 254869 612 254897
rect 646 254869 674 254897
rect 708 254869 736 254897
rect 522 254807 550 254835
rect 584 254807 612 254835
rect 646 254807 674 254835
rect 708 254807 736 254835
rect 522 254745 550 254773
rect 584 254745 612 254773
rect 646 254745 674 254773
rect 708 254745 736 254773
rect 522 245931 550 245959
rect 584 245931 612 245959
rect 646 245931 674 245959
rect 708 245931 736 245959
rect 522 245869 550 245897
rect 584 245869 612 245897
rect 646 245869 674 245897
rect 708 245869 736 245897
rect 522 245807 550 245835
rect 584 245807 612 245835
rect 646 245807 674 245835
rect 708 245807 736 245835
rect 522 245745 550 245773
rect 584 245745 612 245773
rect 646 245745 674 245773
rect 708 245745 736 245773
rect 522 236931 550 236959
rect 584 236931 612 236959
rect 646 236931 674 236959
rect 708 236931 736 236959
rect 522 236869 550 236897
rect 584 236869 612 236897
rect 646 236869 674 236897
rect 708 236869 736 236897
rect 522 236807 550 236835
rect 584 236807 612 236835
rect 646 236807 674 236835
rect 708 236807 736 236835
rect 522 236745 550 236773
rect 584 236745 612 236773
rect 646 236745 674 236773
rect 708 236745 736 236773
rect 522 227931 550 227959
rect 584 227931 612 227959
rect 646 227931 674 227959
rect 708 227931 736 227959
rect 522 227869 550 227897
rect 584 227869 612 227897
rect 646 227869 674 227897
rect 708 227869 736 227897
rect 522 227807 550 227835
rect 584 227807 612 227835
rect 646 227807 674 227835
rect 708 227807 736 227835
rect 522 227745 550 227773
rect 584 227745 612 227773
rect 646 227745 674 227773
rect 708 227745 736 227773
rect 522 218931 550 218959
rect 584 218931 612 218959
rect 646 218931 674 218959
rect 708 218931 736 218959
rect 522 218869 550 218897
rect 584 218869 612 218897
rect 646 218869 674 218897
rect 708 218869 736 218897
rect 522 218807 550 218835
rect 584 218807 612 218835
rect 646 218807 674 218835
rect 708 218807 736 218835
rect 522 218745 550 218773
rect 584 218745 612 218773
rect 646 218745 674 218773
rect 708 218745 736 218773
rect 522 209931 550 209959
rect 584 209931 612 209959
rect 646 209931 674 209959
rect 708 209931 736 209959
rect 522 209869 550 209897
rect 584 209869 612 209897
rect 646 209869 674 209897
rect 708 209869 736 209897
rect 522 209807 550 209835
rect 584 209807 612 209835
rect 646 209807 674 209835
rect 708 209807 736 209835
rect 522 209745 550 209773
rect 584 209745 612 209773
rect 646 209745 674 209773
rect 708 209745 736 209773
rect 522 200931 550 200959
rect 584 200931 612 200959
rect 646 200931 674 200959
rect 708 200931 736 200959
rect 522 200869 550 200897
rect 584 200869 612 200897
rect 646 200869 674 200897
rect 708 200869 736 200897
rect 522 200807 550 200835
rect 584 200807 612 200835
rect 646 200807 674 200835
rect 708 200807 736 200835
rect 522 200745 550 200773
rect 584 200745 612 200773
rect 646 200745 674 200773
rect 708 200745 736 200773
rect 522 191931 550 191959
rect 584 191931 612 191959
rect 646 191931 674 191959
rect 708 191931 736 191959
rect 522 191869 550 191897
rect 584 191869 612 191897
rect 646 191869 674 191897
rect 708 191869 736 191897
rect 522 191807 550 191835
rect 584 191807 612 191835
rect 646 191807 674 191835
rect 708 191807 736 191835
rect 522 191745 550 191773
rect 584 191745 612 191773
rect 646 191745 674 191773
rect 708 191745 736 191773
rect 522 182931 550 182959
rect 584 182931 612 182959
rect 646 182931 674 182959
rect 708 182931 736 182959
rect 522 182869 550 182897
rect 584 182869 612 182897
rect 646 182869 674 182897
rect 708 182869 736 182897
rect 522 182807 550 182835
rect 584 182807 612 182835
rect 646 182807 674 182835
rect 708 182807 736 182835
rect 522 182745 550 182773
rect 584 182745 612 182773
rect 646 182745 674 182773
rect 708 182745 736 182773
rect 522 173931 550 173959
rect 584 173931 612 173959
rect 646 173931 674 173959
rect 708 173931 736 173959
rect 522 173869 550 173897
rect 584 173869 612 173897
rect 646 173869 674 173897
rect 708 173869 736 173897
rect 522 173807 550 173835
rect 584 173807 612 173835
rect 646 173807 674 173835
rect 708 173807 736 173835
rect 522 173745 550 173773
rect 584 173745 612 173773
rect 646 173745 674 173773
rect 708 173745 736 173773
rect 522 164931 550 164959
rect 584 164931 612 164959
rect 646 164931 674 164959
rect 708 164931 736 164959
rect 522 164869 550 164897
rect 584 164869 612 164897
rect 646 164869 674 164897
rect 708 164869 736 164897
rect 522 164807 550 164835
rect 584 164807 612 164835
rect 646 164807 674 164835
rect 708 164807 736 164835
rect 522 164745 550 164773
rect 584 164745 612 164773
rect 646 164745 674 164773
rect 708 164745 736 164773
rect 522 155931 550 155959
rect 584 155931 612 155959
rect 646 155931 674 155959
rect 708 155931 736 155959
rect 522 155869 550 155897
rect 584 155869 612 155897
rect 646 155869 674 155897
rect 708 155869 736 155897
rect 522 155807 550 155835
rect 584 155807 612 155835
rect 646 155807 674 155835
rect 708 155807 736 155835
rect 522 155745 550 155773
rect 584 155745 612 155773
rect 646 155745 674 155773
rect 708 155745 736 155773
rect 522 146931 550 146959
rect 584 146931 612 146959
rect 646 146931 674 146959
rect 708 146931 736 146959
rect 522 146869 550 146897
rect 584 146869 612 146897
rect 646 146869 674 146897
rect 708 146869 736 146897
rect 522 146807 550 146835
rect 584 146807 612 146835
rect 646 146807 674 146835
rect 708 146807 736 146835
rect 522 146745 550 146773
rect 584 146745 612 146773
rect 646 146745 674 146773
rect 708 146745 736 146773
rect 522 137931 550 137959
rect 584 137931 612 137959
rect 646 137931 674 137959
rect 708 137931 736 137959
rect 522 137869 550 137897
rect 584 137869 612 137897
rect 646 137869 674 137897
rect 708 137869 736 137897
rect 522 137807 550 137835
rect 584 137807 612 137835
rect 646 137807 674 137835
rect 708 137807 736 137835
rect 522 137745 550 137773
rect 584 137745 612 137773
rect 646 137745 674 137773
rect 708 137745 736 137773
rect 522 128931 550 128959
rect 584 128931 612 128959
rect 646 128931 674 128959
rect 708 128931 736 128959
rect 522 128869 550 128897
rect 584 128869 612 128897
rect 646 128869 674 128897
rect 708 128869 736 128897
rect 522 128807 550 128835
rect 584 128807 612 128835
rect 646 128807 674 128835
rect 708 128807 736 128835
rect 522 128745 550 128773
rect 584 128745 612 128773
rect 646 128745 674 128773
rect 708 128745 736 128773
rect 522 119931 550 119959
rect 584 119931 612 119959
rect 646 119931 674 119959
rect 708 119931 736 119959
rect 522 119869 550 119897
rect 584 119869 612 119897
rect 646 119869 674 119897
rect 708 119869 736 119897
rect 522 119807 550 119835
rect 584 119807 612 119835
rect 646 119807 674 119835
rect 708 119807 736 119835
rect 522 119745 550 119773
rect 584 119745 612 119773
rect 646 119745 674 119773
rect 708 119745 736 119773
rect 522 110931 550 110959
rect 584 110931 612 110959
rect 646 110931 674 110959
rect 708 110931 736 110959
rect 522 110869 550 110897
rect 584 110869 612 110897
rect 646 110869 674 110897
rect 708 110869 736 110897
rect 522 110807 550 110835
rect 584 110807 612 110835
rect 646 110807 674 110835
rect 708 110807 736 110835
rect 522 110745 550 110773
rect 584 110745 612 110773
rect 646 110745 674 110773
rect 708 110745 736 110773
rect 522 101931 550 101959
rect 584 101931 612 101959
rect 646 101931 674 101959
rect 708 101931 736 101959
rect 522 101869 550 101897
rect 584 101869 612 101897
rect 646 101869 674 101897
rect 708 101869 736 101897
rect 522 101807 550 101835
rect 584 101807 612 101835
rect 646 101807 674 101835
rect 708 101807 736 101835
rect 522 101745 550 101773
rect 584 101745 612 101773
rect 646 101745 674 101773
rect 708 101745 736 101773
rect 522 92931 550 92959
rect 584 92931 612 92959
rect 646 92931 674 92959
rect 708 92931 736 92959
rect 522 92869 550 92897
rect 584 92869 612 92897
rect 646 92869 674 92897
rect 708 92869 736 92897
rect 522 92807 550 92835
rect 584 92807 612 92835
rect 646 92807 674 92835
rect 708 92807 736 92835
rect 522 92745 550 92773
rect 584 92745 612 92773
rect 646 92745 674 92773
rect 708 92745 736 92773
rect 522 83931 550 83959
rect 584 83931 612 83959
rect 646 83931 674 83959
rect 708 83931 736 83959
rect 522 83869 550 83897
rect 584 83869 612 83897
rect 646 83869 674 83897
rect 708 83869 736 83897
rect 522 83807 550 83835
rect 584 83807 612 83835
rect 646 83807 674 83835
rect 708 83807 736 83835
rect 522 83745 550 83773
rect 584 83745 612 83773
rect 646 83745 674 83773
rect 708 83745 736 83773
rect 522 74931 550 74959
rect 584 74931 612 74959
rect 646 74931 674 74959
rect 708 74931 736 74959
rect 522 74869 550 74897
rect 584 74869 612 74897
rect 646 74869 674 74897
rect 708 74869 736 74897
rect 522 74807 550 74835
rect 584 74807 612 74835
rect 646 74807 674 74835
rect 708 74807 736 74835
rect 522 74745 550 74773
rect 584 74745 612 74773
rect 646 74745 674 74773
rect 708 74745 736 74773
rect 522 65931 550 65959
rect 584 65931 612 65959
rect 646 65931 674 65959
rect 708 65931 736 65959
rect 522 65869 550 65897
rect 584 65869 612 65897
rect 646 65869 674 65897
rect 708 65869 736 65897
rect 522 65807 550 65835
rect 584 65807 612 65835
rect 646 65807 674 65835
rect 708 65807 736 65835
rect 522 65745 550 65773
rect 584 65745 612 65773
rect 646 65745 674 65773
rect 708 65745 736 65773
rect 522 56931 550 56959
rect 584 56931 612 56959
rect 646 56931 674 56959
rect 708 56931 736 56959
rect 522 56869 550 56897
rect 584 56869 612 56897
rect 646 56869 674 56897
rect 708 56869 736 56897
rect 522 56807 550 56835
rect 584 56807 612 56835
rect 646 56807 674 56835
rect 708 56807 736 56835
rect 522 56745 550 56773
rect 584 56745 612 56773
rect 646 56745 674 56773
rect 708 56745 736 56773
rect 522 47931 550 47959
rect 584 47931 612 47959
rect 646 47931 674 47959
rect 708 47931 736 47959
rect 522 47869 550 47897
rect 584 47869 612 47897
rect 646 47869 674 47897
rect 708 47869 736 47897
rect 522 47807 550 47835
rect 584 47807 612 47835
rect 646 47807 674 47835
rect 708 47807 736 47835
rect 522 47745 550 47773
rect 584 47745 612 47773
rect 646 47745 674 47773
rect 708 47745 736 47773
rect 522 38931 550 38959
rect 584 38931 612 38959
rect 646 38931 674 38959
rect 708 38931 736 38959
rect 522 38869 550 38897
rect 584 38869 612 38897
rect 646 38869 674 38897
rect 708 38869 736 38897
rect 522 38807 550 38835
rect 584 38807 612 38835
rect 646 38807 674 38835
rect 708 38807 736 38835
rect 522 38745 550 38773
rect 584 38745 612 38773
rect 646 38745 674 38773
rect 708 38745 736 38773
rect 522 29931 550 29959
rect 584 29931 612 29959
rect 646 29931 674 29959
rect 708 29931 736 29959
rect 522 29869 550 29897
rect 584 29869 612 29897
rect 646 29869 674 29897
rect 708 29869 736 29897
rect 522 29807 550 29835
rect 584 29807 612 29835
rect 646 29807 674 29835
rect 708 29807 736 29835
rect 522 29745 550 29773
rect 584 29745 612 29773
rect 646 29745 674 29773
rect 708 29745 736 29773
rect 522 20931 550 20959
rect 584 20931 612 20959
rect 646 20931 674 20959
rect 708 20931 736 20959
rect 522 20869 550 20897
rect 584 20869 612 20897
rect 646 20869 674 20897
rect 708 20869 736 20897
rect 522 20807 550 20835
rect 584 20807 612 20835
rect 646 20807 674 20835
rect 708 20807 736 20835
rect 522 20745 550 20773
rect 584 20745 612 20773
rect 646 20745 674 20773
rect 708 20745 736 20773
rect 522 11931 550 11959
rect 584 11931 612 11959
rect 646 11931 674 11959
rect 708 11931 736 11959
rect 522 11869 550 11897
rect 584 11869 612 11897
rect 646 11869 674 11897
rect 708 11869 736 11897
rect 522 11807 550 11835
rect 584 11807 612 11835
rect 646 11807 674 11835
rect 708 11807 736 11835
rect 522 11745 550 11773
rect 584 11745 612 11773
rect 646 11745 674 11773
rect 708 11745 736 11773
rect 522 2931 550 2959
rect 584 2931 612 2959
rect 646 2931 674 2959
rect 708 2931 736 2959
rect 522 2869 550 2897
rect 584 2869 612 2897
rect 646 2869 674 2897
rect 708 2869 736 2897
rect 522 2807 550 2835
rect 584 2807 612 2835
rect 646 2807 674 2835
rect 708 2807 736 2835
rect 522 2745 550 2773
rect 584 2745 612 2773
rect 646 2745 674 2773
rect 708 2745 736 2773
rect 522 876 550 904
rect 584 876 612 904
rect 646 876 674 904
rect 708 876 736 904
rect 522 814 550 842
rect 584 814 612 842
rect 646 814 674 842
rect 708 814 736 842
rect 522 752 550 780
rect 584 752 612 780
rect 646 752 674 780
rect 708 752 736 780
rect 522 690 550 718
rect 584 690 612 718
rect 646 690 674 718
rect 708 690 736 718
rect 2577 299162 2605 299190
rect 2639 299162 2667 299190
rect 2701 299162 2729 299190
rect 2763 299162 2791 299190
rect 2577 299100 2605 299128
rect 2639 299100 2667 299128
rect 2701 299100 2729 299128
rect 2763 299100 2791 299128
rect 2577 299038 2605 299066
rect 2639 299038 2667 299066
rect 2701 299038 2729 299066
rect 2763 299038 2791 299066
rect 2577 298976 2605 299004
rect 2639 298976 2667 299004
rect 2701 298976 2729 299004
rect 2763 298976 2791 299004
rect 2577 290931 2605 290959
rect 2639 290931 2667 290959
rect 2701 290931 2729 290959
rect 2763 290931 2791 290959
rect 2577 290869 2605 290897
rect 2639 290869 2667 290897
rect 2701 290869 2729 290897
rect 2763 290869 2791 290897
rect 2577 290807 2605 290835
rect 2639 290807 2667 290835
rect 2701 290807 2729 290835
rect 2763 290807 2791 290835
rect 2577 290745 2605 290773
rect 2639 290745 2667 290773
rect 2701 290745 2729 290773
rect 2763 290745 2791 290773
rect 2577 281931 2605 281959
rect 2639 281931 2667 281959
rect 2701 281931 2729 281959
rect 2763 281931 2791 281959
rect 2577 281869 2605 281897
rect 2639 281869 2667 281897
rect 2701 281869 2729 281897
rect 2763 281869 2791 281897
rect 2577 281807 2605 281835
rect 2639 281807 2667 281835
rect 2701 281807 2729 281835
rect 2763 281807 2791 281835
rect 2577 281745 2605 281773
rect 2639 281745 2667 281773
rect 2701 281745 2729 281773
rect 2763 281745 2791 281773
rect 2577 272931 2605 272959
rect 2639 272931 2667 272959
rect 2701 272931 2729 272959
rect 2763 272931 2791 272959
rect 2577 272869 2605 272897
rect 2639 272869 2667 272897
rect 2701 272869 2729 272897
rect 2763 272869 2791 272897
rect 2577 272807 2605 272835
rect 2639 272807 2667 272835
rect 2701 272807 2729 272835
rect 2763 272807 2791 272835
rect 2577 272745 2605 272773
rect 2639 272745 2667 272773
rect 2701 272745 2729 272773
rect 2763 272745 2791 272773
rect 2577 263931 2605 263959
rect 2639 263931 2667 263959
rect 2701 263931 2729 263959
rect 2763 263931 2791 263959
rect 2577 263869 2605 263897
rect 2639 263869 2667 263897
rect 2701 263869 2729 263897
rect 2763 263869 2791 263897
rect 2577 263807 2605 263835
rect 2639 263807 2667 263835
rect 2701 263807 2729 263835
rect 2763 263807 2791 263835
rect 2577 263745 2605 263773
rect 2639 263745 2667 263773
rect 2701 263745 2729 263773
rect 2763 263745 2791 263773
rect 2577 254931 2605 254959
rect 2639 254931 2667 254959
rect 2701 254931 2729 254959
rect 2763 254931 2791 254959
rect 2577 254869 2605 254897
rect 2639 254869 2667 254897
rect 2701 254869 2729 254897
rect 2763 254869 2791 254897
rect 2577 254807 2605 254835
rect 2639 254807 2667 254835
rect 2701 254807 2729 254835
rect 2763 254807 2791 254835
rect 2577 254745 2605 254773
rect 2639 254745 2667 254773
rect 2701 254745 2729 254773
rect 2763 254745 2791 254773
rect 2577 245931 2605 245959
rect 2639 245931 2667 245959
rect 2701 245931 2729 245959
rect 2763 245931 2791 245959
rect 2577 245869 2605 245897
rect 2639 245869 2667 245897
rect 2701 245869 2729 245897
rect 2763 245869 2791 245897
rect 2577 245807 2605 245835
rect 2639 245807 2667 245835
rect 2701 245807 2729 245835
rect 2763 245807 2791 245835
rect 2577 245745 2605 245773
rect 2639 245745 2667 245773
rect 2701 245745 2729 245773
rect 2763 245745 2791 245773
rect 2577 236931 2605 236959
rect 2639 236931 2667 236959
rect 2701 236931 2729 236959
rect 2763 236931 2791 236959
rect 2577 236869 2605 236897
rect 2639 236869 2667 236897
rect 2701 236869 2729 236897
rect 2763 236869 2791 236897
rect 2577 236807 2605 236835
rect 2639 236807 2667 236835
rect 2701 236807 2729 236835
rect 2763 236807 2791 236835
rect 2577 236745 2605 236773
rect 2639 236745 2667 236773
rect 2701 236745 2729 236773
rect 2763 236745 2791 236773
rect 2577 227931 2605 227959
rect 2639 227931 2667 227959
rect 2701 227931 2729 227959
rect 2763 227931 2791 227959
rect 2577 227869 2605 227897
rect 2639 227869 2667 227897
rect 2701 227869 2729 227897
rect 2763 227869 2791 227897
rect 2577 227807 2605 227835
rect 2639 227807 2667 227835
rect 2701 227807 2729 227835
rect 2763 227807 2791 227835
rect 2577 227745 2605 227773
rect 2639 227745 2667 227773
rect 2701 227745 2729 227773
rect 2763 227745 2791 227773
rect 2577 218931 2605 218959
rect 2639 218931 2667 218959
rect 2701 218931 2729 218959
rect 2763 218931 2791 218959
rect 2577 218869 2605 218897
rect 2639 218869 2667 218897
rect 2701 218869 2729 218897
rect 2763 218869 2791 218897
rect 2577 218807 2605 218835
rect 2639 218807 2667 218835
rect 2701 218807 2729 218835
rect 2763 218807 2791 218835
rect 2577 218745 2605 218773
rect 2639 218745 2667 218773
rect 2701 218745 2729 218773
rect 2763 218745 2791 218773
rect 2577 209931 2605 209959
rect 2639 209931 2667 209959
rect 2701 209931 2729 209959
rect 2763 209931 2791 209959
rect 2577 209869 2605 209897
rect 2639 209869 2667 209897
rect 2701 209869 2729 209897
rect 2763 209869 2791 209897
rect 2577 209807 2605 209835
rect 2639 209807 2667 209835
rect 2701 209807 2729 209835
rect 2763 209807 2791 209835
rect 2577 209745 2605 209773
rect 2639 209745 2667 209773
rect 2701 209745 2729 209773
rect 2763 209745 2791 209773
rect 2577 200931 2605 200959
rect 2639 200931 2667 200959
rect 2701 200931 2729 200959
rect 2763 200931 2791 200959
rect 2577 200869 2605 200897
rect 2639 200869 2667 200897
rect 2701 200869 2729 200897
rect 2763 200869 2791 200897
rect 2577 200807 2605 200835
rect 2639 200807 2667 200835
rect 2701 200807 2729 200835
rect 2763 200807 2791 200835
rect 2577 200745 2605 200773
rect 2639 200745 2667 200773
rect 2701 200745 2729 200773
rect 2763 200745 2791 200773
rect 2577 191931 2605 191959
rect 2639 191931 2667 191959
rect 2701 191931 2729 191959
rect 2763 191931 2791 191959
rect 2577 191869 2605 191897
rect 2639 191869 2667 191897
rect 2701 191869 2729 191897
rect 2763 191869 2791 191897
rect 2577 191807 2605 191835
rect 2639 191807 2667 191835
rect 2701 191807 2729 191835
rect 2763 191807 2791 191835
rect 2577 191745 2605 191773
rect 2639 191745 2667 191773
rect 2701 191745 2729 191773
rect 2763 191745 2791 191773
rect 2577 182931 2605 182959
rect 2639 182931 2667 182959
rect 2701 182931 2729 182959
rect 2763 182931 2791 182959
rect 2577 182869 2605 182897
rect 2639 182869 2667 182897
rect 2701 182869 2729 182897
rect 2763 182869 2791 182897
rect 2577 182807 2605 182835
rect 2639 182807 2667 182835
rect 2701 182807 2729 182835
rect 2763 182807 2791 182835
rect 2577 182745 2605 182773
rect 2639 182745 2667 182773
rect 2701 182745 2729 182773
rect 2763 182745 2791 182773
rect 2577 173931 2605 173959
rect 2639 173931 2667 173959
rect 2701 173931 2729 173959
rect 2763 173931 2791 173959
rect 2577 173869 2605 173897
rect 2639 173869 2667 173897
rect 2701 173869 2729 173897
rect 2763 173869 2791 173897
rect 2577 173807 2605 173835
rect 2639 173807 2667 173835
rect 2701 173807 2729 173835
rect 2763 173807 2791 173835
rect 2577 173745 2605 173773
rect 2639 173745 2667 173773
rect 2701 173745 2729 173773
rect 2763 173745 2791 173773
rect 2577 164931 2605 164959
rect 2639 164931 2667 164959
rect 2701 164931 2729 164959
rect 2763 164931 2791 164959
rect 2577 164869 2605 164897
rect 2639 164869 2667 164897
rect 2701 164869 2729 164897
rect 2763 164869 2791 164897
rect 2577 164807 2605 164835
rect 2639 164807 2667 164835
rect 2701 164807 2729 164835
rect 2763 164807 2791 164835
rect 2577 164745 2605 164773
rect 2639 164745 2667 164773
rect 2701 164745 2729 164773
rect 2763 164745 2791 164773
rect 2577 155931 2605 155959
rect 2639 155931 2667 155959
rect 2701 155931 2729 155959
rect 2763 155931 2791 155959
rect 2577 155869 2605 155897
rect 2639 155869 2667 155897
rect 2701 155869 2729 155897
rect 2763 155869 2791 155897
rect 2577 155807 2605 155835
rect 2639 155807 2667 155835
rect 2701 155807 2729 155835
rect 2763 155807 2791 155835
rect 2577 155745 2605 155773
rect 2639 155745 2667 155773
rect 2701 155745 2729 155773
rect 2763 155745 2791 155773
rect 2577 146931 2605 146959
rect 2639 146931 2667 146959
rect 2701 146931 2729 146959
rect 2763 146931 2791 146959
rect 2577 146869 2605 146897
rect 2639 146869 2667 146897
rect 2701 146869 2729 146897
rect 2763 146869 2791 146897
rect 2577 146807 2605 146835
rect 2639 146807 2667 146835
rect 2701 146807 2729 146835
rect 2763 146807 2791 146835
rect 2577 146745 2605 146773
rect 2639 146745 2667 146773
rect 2701 146745 2729 146773
rect 2763 146745 2791 146773
rect 2577 137931 2605 137959
rect 2639 137931 2667 137959
rect 2701 137931 2729 137959
rect 2763 137931 2791 137959
rect 2577 137869 2605 137897
rect 2639 137869 2667 137897
rect 2701 137869 2729 137897
rect 2763 137869 2791 137897
rect 2577 137807 2605 137835
rect 2639 137807 2667 137835
rect 2701 137807 2729 137835
rect 2763 137807 2791 137835
rect 2577 137745 2605 137773
rect 2639 137745 2667 137773
rect 2701 137745 2729 137773
rect 2763 137745 2791 137773
rect 2577 128931 2605 128959
rect 2639 128931 2667 128959
rect 2701 128931 2729 128959
rect 2763 128931 2791 128959
rect 2577 128869 2605 128897
rect 2639 128869 2667 128897
rect 2701 128869 2729 128897
rect 2763 128869 2791 128897
rect 2577 128807 2605 128835
rect 2639 128807 2667 128835
rect 2701 128807 2729 128835
rect 2763 128807 2791 128835
rect 2577 128745 2605 128773
rect 2639 128745 2667 128773
rect 2701 128745 2729 128773
rect 2763 128745 2791 128773
rect 2577 119931 2605 119959
rect 2639 119931 2667 119959
rect 2701 119931 2729 119959
rect 2763 119931 2791 119959
rect 2577 119869 2605 119897
rect 2639 119869 2667 119897
rect 2701 119869 2729 119897
rect 2763 119869 2791 119897
rect 2577 119807 2605 119835
rect 2639 119807 2667 119835
rect 2701 119807 2729 119835
rect 2763 119807 2791 119835
rect 2577 119745 2605 119773
rect 2639 119745 2667 119773
rect 2701 119745 2729 119773
rect 2763 119745 2791 119773
rect 2577 110931 2605 110959
rect 2639 110931 2667 110959
rect 2701 110931 2729 110959
rect 2763 110931 2791 110959
rect 2577 110869 2605 110897
rect 2639 110869 2667 110897
rect 2701 110869 2729 110897
rect 2763 110869 2791 110897
rect 2577 110807 2605 110835
rect 2639 110807 2667 110835
rect 2701 110807 2729 110835
rect 2763 110807 2791 110835
rect 2577 110745 2605 110773
rect 2639 110745 2667 110773
rect 2701 110745 2729 110773
rect 2763 110745 2791 110773
rect 2577 101931 2605 101959
rect 2639 101931 2667 101959
rect 2701 101931 2729 101959
rect 2763 101931 2791 101959
rect 2577 101869 2605 101897
rect 2639 101869 2667 101897
rect 2701 101869 2729 101897
rect 2763 101869 2791 101897
rect 2577 101807 2605 101835
rect 2639 101807 2667 101835
rect 2701 101807 2729 101835
rect 2763 101807 2791 101835
rect 2577 101745 2605 101773
rect 2639 101745 2667 101773
rect 2701 101745 2729 101773
rect 2763 101745 2791 101773
rect 2577 92931 2605 92959
rect 2639 92931 2667 92959
rect 2701 92931 2729 92959
rect 2763 92931 2791 92959
rect 2577 92869 2605 92897
rect 2639 92869 2667 92897
rect 2701 92869 2729 92897
rect 2763 92869 2791 92897
rect 2577 92807 2605 92835
rect 2639 92807 2667 92835
rect 2701 92807 2729 92835
rect 2763 92807 2791 92835
rect 2577 92745 2605 92773
rect 2639 92745 2667 92773
rect 2701 92745 2729 92773
rect 2763 92745 2791 92773
rect 2577 83931 2605 83959
rect 2639 83931 2667 83959
rect 2701 83931 2729 83959
rect 2763 83931 2791 83959
rect 2577 83869 2605 83897
rect 2639 83869 2667 83897
rect 2701 83869 2729 83897
rect 2763 83869 2791 83897
rect 2577 83807 2605 83835
rect 2639 83807 2667 83835
rect 2701 83807 2729 83835
rect 2763 83807 2791 83835
rect 2577 83745 2605 83773
rect 2639 83745 2667 83773
rect 2701 83745 2729 83773
rect 2763 83745 2791 83773
rect 2577 74931 2605 74959
rect 2639 74931 2667 74959
rect 2701 74931 2729 74959
rect 2763 74931 2791 74959
rect 2577 74869 2605 74897
rect 2639 74869 2667 74897
rect 2701 74869 2729 74897
rect 2763 74869 2791 74897
rect 2577 74807 2605 74835
rect 2639 74807 2667 74835
rect 2701 74807 2729 74835
rect 2763 74807 2791 74835
rect 2577 74745 2605 74773
rect 2639 74745 2667 74773
rect 2701 74745 2729 74773
rect 2763 74745 2791 74773
rect 2577 65931 2605 65959
rect 2639 65931 2667 65959
rect 2701 65931 2729 65959
rect 2763 65931 2791 65959
rect 2577 65869 2605 65897
rect 2639 65869 2667 65897
rect 2701 65869 2729 65897
rect 2763 65869 2791 65897
rect 2577 65807 2605 65835
rect 2639 65807 2667 65835
rect 2701 65807 2729 65835
rect 2763 65807 2791 65835
rect 2577 65745 2605 65773
rect 2639 65745 2667 65773
rect 2701 65745 2729 65773
rect 2763 65745 2791 65773
rect 2577 56931 2605 56959
rect 2639 56931 2667 56959
rect 2701 56931 2729 56959
rect 2763 56931 2791 56959
rect 2577 56869 2605 56897
rect 2639 56869 2667 56897
rect 2701 56869 2729 56897
rect 2763 56869 2791 56897
rect 2577 56807 2605 56835
rect 2639 56807 2667 56835
rect 2701 56807 2729 56835
rect 2763 56807 2791 56835
rect 2577 56745 2605 56773
rect 2639 56745 2667 56773
rect 2701 56745 2729 56773
rect 2763 56745 2791 56773
rect 2577 47931 2605 47959
rect 2639 47931 2667 47959
rect 2701 47931 2729 47959
rect 2763 47931 2791 47959
rect 2577 47869 2605 47897
rect 2639 47869 2667 47897
rect 2701 47869 2729 47897
rect 2763 47869 2791 47897
rect 2577 47807 2605 47835
rect 2639 47807 2667 47835
rect 2701 47807 2729 47835
rect 2763 47807 2791 47835
rect 2577 47745 2605 47773
rect 2639 47745 2667 47773
rect 2701 47745 2729 47773
rect 2763 47745 2791 47773
rect 2577 38931 2605 38959
rect 2639 38931 2667 38959
rect 2701 38931 2729 38959
rect 2763 38931 2791 38959
rect 2577 38869 2605 38897
rect 2639 38869 2667 38897
rect 2701 38869 2729 38897
rect 2763 38869 2791 38897
rect 2577 38807 2605 38835
rect 2639 38807 2667 38835
rect 2701 38807 2729 38835
rect 2763 38807 2791 38835
rect 2577 38745 2605 38773
rect 2639 38745 2667 38773
rect 2701 38745 2729 38773
rect 2763 38745 2791 38773
rect 2577 29931 2605 29959
rect 2639 29931 2667 29959
rect 2701 29931 2729 29959
rect 2763 29931 2791 29959
rect 2577 29869 2605 29897
rect 2639 29869 2667 29897
rect 2701 29869 2729 29897
rect 2763 29869 2791 29897
rect 2577 29807 2605 29835
rect 2639 29807 2667 29835
rect 2701 29807 2729 29835
rect 2763 29807 2791 29835
rect 2577 29745 2605 29773
rect 2639 29745 2667 29773
rect 2701 29745 2729 29773
rect 2763 29745 2791 29773
rect 2577 20931 2605 20959
rect 2639 20931 2667 20959
rect 2701 20931 2729 20959
rect 2763 20931 2791 20959
rect 2577 20869 2605 20897
rect 2639 20869 2667 20897
rect 2701 20869 2729 20897
rect 2763 20869 2791 20897
rect 2577 20807 2605 20835
rect 2639 20807 2667 20835
rect 2701 20807 2729 20835
rect 2763 20807 2791 20835
rect 2577 20745 2605 20773
rect 2639 20745 2667 20773
rect 2701 20745 2729 20773
rect 2763 20745 2791 20773
rect 2577 11931 2605 11959
rect 2639 11931 2667 11959
rect 2701 11931 2729 11959
rect 2763 11931 2791 11959
rect 2577 11869 2605 11897
rect 2639 11869 2667 11897
rect 2701 11869 2729 11897
rect 2763 11869 2791 11897
rect 2577 11807 2605 11835
rect 2639 11807 2667 11835
rect 2701 11807 2729 11835
rect 2763 11807 2791 11835
rect 2577 11745 2605 11773
rect 2639 11745 2667 11773
rect 2701 11745 2729 11773
rect 2763 11745 2791 11773
rect 2577 2931 2605 2959
rect 2639 2931 2667 2959
rect 2701 2931 2729 2959
rect 2763 2931 2791 2959
rect 2577 2869 2605 2897
rect 2639 2869 2667 2897
rect 2701 2869 2729 2897
rect 2763 2869 2791 2897
rect 2577 2807 2605 2835
rect 2639 2807 2667 2835
rect 2701 2807 2729 2835
rect 2763 2807 2791 2835
rect 2577 2745 2605 2773
rect 2639 2745 2667 2773
rect 2701 2745 2729 2773
rect 2763 2745 2791 2773
rect 2577 876 2605 904
rect 2639 876 2667 904
rect 2701 876 2729 904
rect 2763 876 2791 904
rect 2577 814 2605 842
rect 2639 814 2667 842
rect 2701 814 2729 842
rect 2763 814 2791 842
rect 2577 752 2605 780
rect 2639 752 2667 780
rect 2701 752 2729 780
rect 2763 752 2791 780
rect 2577 690 2605 718
rect 2639 690 2667 718
rect 2701 690 2729 718
rect 2763 690 2791 718
rect 42 396 70 424
rect 104 396 132 424
rect 166 396 194 424
rect 228 396 256 424
rect 42 334 70 362
rect 104 334 132 362
rect 166 334 194 362
rect 228 334 256 362
rect 42 272 70 300
rect 104 272 132 300
rect 166 272 194 300
rect 228 272 256 300
rect 42 210 70 238
rect 104 210 132 238
rect 166 210 194 238
rect 228 210 256 238
rect 4437 299642 4465 299670
rect 4499 299642 4527 299670
rect 4561 299642 4589 299670
rect 4623 299642 4651 299670
rect 4437 299580 4465 299608
rect 4499 299580 4527 299608
rect 4561 299580 4589 299608
rect 4623 299580 4651 299608
rect 4437 299518 4465 299546
rect 4499 299518 4527 299546
rect 4561 299518 4589 299546
rect 4623 299518 4651 299546
rect 4437 299456 4465 299484
rect 4499 299456 4527 299484
rect 4561 299456 4589 299484
rect 4623 299456 4651 299484
rect 4437 293931 4465 293959
rect 4499 293931 4527 293959
rect 4561 293931 4589 293959
rect 4623 293931 4651 293959
rect 4437 293869 4465 293897
rect 4499 293869 4527 293897
rect 4561 293869 4589 293897
rect 4623 293869 4651 293897
rect 4437 293807 4465 293835
rect 4499 293807 4527 293835
rect 4561 293807 4589 293835
rect 4623 293807 4651 293835
rect 4437 293745 4465 293773
rect 4499 293745 4527 293773
rect 4561 293745 4589 293773
rect 4623 293745 4651 293773
rect 4437 284931 4465 284959
rect 4499 284931 4527 284959
rect 4561 284931 4589 284959
rect 4623 284931 4651 284959
rect 4437 284869 4465 284897
rect 4499 284869 4527 284897
rect 4561 284869 4589 284897
rect 4623 284869 4651 284897
rect 4437 284807 4465 284835
rect 4499 284807 4527 284835
rect 4561 284807 4589 284835
rect 4623 284807 4651 284835
rect 4437 284745 4465 284773
rect 4499 284745 4527 284773
rect 4561 284745 4589 284773
rect 4623 284745 4651 284773
rect 4437 275931 4465 275959
rect 4499 275931 4527 275959
rect 4561 275931 4589 275959
rect 4623 275931 4651 275959
rect 4437 275869 4465 275897
rect 4499 275869 4527 275897
rect 4561 275869 4589 275897
rect 4623 275869 4651 275897
rect 4437 275807 4465 275835
rect 4499 275807 4527 275835
rect 4561 275807 4589 275835
rect 4623 275807 4651 275835
rect 4437 275745 4465 275773
rect 4499 275745 4527 275773
rect 4561 275745 4589 275773
rect 4623 275745 4651 275773
rect 4437 266931 4465 266959
rect 4499 266931 4527 266959
rect 4561 266931 4589 266959
rect 4623 266931 4651 266959
rect 4437 266869 4465 266897
rect 4499 266869 4527 266897
rect 4561 266869 4589 266897
rect 4623 266869 4651 266897
rect 4437 266807 4465 266835
rect 4499 266807 4527 266835
rect 4561 266807 4589 266835
rect 4623 266807 4651 266835
rect 4437 266745 4465 266773
rect 4499 266745 4527 266773
rect 4561 266745 4589 266773
rect 4623 266745 4651 266773
rect 4437 257931 4465 257959
rect 4499 257931 4527 257959
rect 4561 257931 4589 257959
rect 4623 257931 4651 257959
rect 4437 257869 4465 257897
rect 4499 257869 4527 257897
rect 4561 257869 4589 257897
rect 4623 257869 4651 257897
rect 4437 257807 4465 257835
rect 4499 257807 4527 257835
rect 4561 257807 4589 257835
rect 4623 257807 4651 257835
rect 4437 257745 4465 257773
rect 4499 257745 4527 257773
rect 4561 257745 4589 257773
rect 4623 257745 4651 257773
rect 4437 248931 4465 248959
rect 4499 248931 4527 248959
rect 4561 248931 4589 248959
rect 4623 248931 4651 248959
rect 4437 248869 4465 248897
rect 4499 248869 4527 248897
rect 4561 248869 4589 248897
rect 4623 248869 4651 248897
rect 4437 248807 4465 248835
rect 4499 248807 4527 248835
rect 4561 248807 4589 248835
rect 4623 248807 4651 248835
rect 4437 248745 4465 248773
rect 4499 248745 4527 248773
rect 4561 248745 4589 248773
rect 4623 248745 4651 248773
rect 4437 239931 4465 239959
rect 4499 239931 4527 239959
rect 4561 239931 4589 239959
rect 4623 239931 4651 239959
rect 4437 239869 4465 239897
rect 4499 239869 4527 239897
rect 4561 239869 4589 239897
rect 4623 239869 4651 239897
rect 4437 239807 4465 239835
rect 4499 239807 4527 239835
rect 4561 239807 4589 239835
rect 4623 239807 4651 239835
rect 4437 239745 4465 239773
rect 4499 239745 4527 239773
rect 4561 239745 4589 239773
rect 4623 239745 4651 239773
rect 4437 230931 4465 230959
rect 4499 230931 4527 230959
rect 4561 230931 4589 230959
rect 4623 230931 4651 230959
rect 4437 230869 4465 230897
rect 4499 230869 4527 230897
rect 4561 230869 4589 230897
rect 4623 230869 4651 230897
rect 4437 230807 4465 230835
rect 4499 230807 4527 230835
rect 4561 230807 4589 230835
rect 4623 230807 4651 230835
rect 4437 230745 4465 230773
rect 4499 230745 4527 230773
rect 4561 230745 4589 230773
rect 4623 230745 4651 230773
rect 4437 221931 4465 221959
rect 4499 221931 4527 221959
rect 4561 221931 4589 221959
rect 4623 221931 4651 221959
rect 4437 221869 4465 221897
rect 4499 221869 4527 221897
rect 4561 221869 4589 221897
rect 4623 221869 4651 221897
rect 4437 221807 4465 221835
rect 4499 221807 4527 221835
rect 4561 221807 4589 221835
rect 4623 221807 4651 221835
rect 4437 221745 4465 221773
rect 4499 221745 4527 221773
rect 4561 221745 4589 221773
rect 4623 221745 4651 221773
rect 4437 212931 4465 212959
rect 4499 212931 4527 212959
rect 4561 212931 4589 212959
rect 4623 212931 4651 212959
rect 4437 212869 4465 212897
rect 4499 212869 4527 212897
rect 4561 212869 4589 212897
rect 4623 212869 4651 212897
rect 4437 212807 4465 212835
rect 4499 212807 4527 212835
rect 4561 212807 4589 212835
rect 4623 212807 4651 212835
rect 4437 212745 4465 212773
rect 4499 212745 4527 212773
rect 4561 212745 4589 212773
rect 4623 212745 4651 212773
rect 4437 203931 4465 203959
rect 4499 203931 4527 203959
rect 4561 203931 4589 203959
rect 4623 203931 4651 203959
rect 4437 203869 4465 203897
rect 4499 203869 4527 203897
rect 4561 203869 4589 203897
rect 4623 203869 4651 203897
rect 4437 203807 4465 203835
rect 4499 203807 4527 203835
rect 4561 203807 4589 203835
rect 4623 203807 4651 203835
rect 4437 203745 4465 203773
rect 4499 203745 4527 203773
rect 4561 203745 4589 203773
rect 4623 203745 4651 203773
rect 4437 194931 4465 194959
rect 4499 194931 4527 194959
rect 4561 194931 4589 194959
rect 4623 194931 4651 194959
rect 4437 194869 4465 194897
rect 4499 194869 4527 194897
rect 4561 194869 4589 194897
rect 4623 194869 4651 194897
rect 4437 194807 4465 194835
rect 4499 194807 4527 194835
rect 4561 194807 4589 194835
rect 4623 194807 4651 194835
rect 4437 194745 4465 194773
rect 4499 194745 4527 194773
rect 4561 194745 4589 194773
rect 4623 194745 4651 194773
rect 4437 185931 4465 185959
rect 4499 185931 4527 185959
rect 4561 185931 4589 185959
rect 4623 185931 4651 185959
rect 4437 185869 4465 185897
rect 4499 185869 4527 185897
rect 4561 185869 4589 185897
rect 4623 185869 4651 185897
rect 4437 185807 4465 185835
rect 4499 185807 4527 185835
rect 4561 185807 4589 185835
rect 4623 185807 4651 185835
rect 4437 185745 4465 185773
rect 4499 185745 4527 185773
rect 4561 185745 4589 185773
rect 4623 185745 4651 185773
rect 4437 176931 4465 176959
rect 4499 176931 4527 176959
rect 4561 176931 4589 176959
rect 4623 176931 4651 176959
rect 4437 176869 4465 176897
rect 4499 176869 4527 176897
rect 4561 176869 4589 176897
rect 4623 176869 4651 176897
rect 4437 176807 4465 176835
rect 4499 176807 4527 176835
rect 4561 176807 4589 176835
rect 4623 176807 4651 176835
rect 4437 176745 4465 176773
rect 4499 176745 4527 176773
rect 4561 176745 4589 176773
rect 4623 176745 4651 176773
rect 4437 167931 4465 167959
rect 4499 167931 4527 167959
rect 4561 167931 4589 167959
rect 4623 167931 4651 167959
rect 4437 167869 4465 167897
rect 4499 167869 4527 167897
rect 4561 167869 4589 167897
rect 4623 167869 4651 167897
rect 4437 167807 4465 167835
rect 4499 167807 4527 167835
rect 4561 167807 4589 167835
rect 4623 167807 4651 167835
rect 4437 167745 4465 167773
rect 4499 167745 4527 167773
rect 4561 167745 4589 167773
rect 4623 167745 4651 167773
rect 4437 158931 4465 158959
rect 4499 158931 4527 158959
rect 4561 158931 4589 158959
rect 4623 158931 4651 158959
rect 4437 158869 4465 158897
rect 4499 158869 4527 158897
rect 4561 158869 4589 158897
rect 4623 158869 4651 158897
rect 4437 158807 4465 158835
rect 4499 158807 4527 158835
rect 4561 158807 4589 158835
rect 4623 158807 4651 158835
rect 4437 158745 4465 158773
rect 4499 158745 4527 158773
rect 4561 158745 4589 158773
rect 4623 158745 4651 158773
rect 4437 149931 4465 149959
rect 4499 149931 4527 149959
rect 4561 149931 4589 149959
rect 4623 149931 4651 149959
rect 4437 149869 4465 149897
rect 4499 149869 4527 149897
rect 4561 149869 4589 149897
rect 4623 149869 4651 149897
rect 4437 149807 4465 149835
rect 4499 149807 4527 149835
rect 4561 149807 4589 149835
rect 4623 149807 4651 149835
rect 4437 149745 4465 149773
rect 4499 149745 4527 149773
rect 4561 149745 4589 149773
rect 4623 149745 4651 149773
rect 4437 140931 4465 140959
rect 4499 140931 4527 140959
rect 4561 140931 4589 140959
rect 4623 140931 4651 140959
rect 4437 140869 4465 140897
rect 4499 140869 4527 140897
rect 4561 140869 4589 140897
rect 4623 140869 4651 140897
rect 4437 140807 4465 140835
rect 4499 140807 4527 140835
rect 4561 140807 4589 140835
rect 4623 140807 4651 140835
rect 4437 140745 4465 140773
rect 4499 140745 4527 140773
rect 4561 140745 4589 140773
rect 4623 140745 4651 140773
rect 4437 131931 4465 131959
rect 4499 131931 4527 131959
rect 4561 131931 4589 131959
rect 4623 131931 4651 131959
rect 4437 131869 4465 131897
rect 4499 131869 4527 131897
rect 4561 131869 4589 131897
rect 4623 131869 4651 131897
rect 4437 131807 4465 131835
rect 4499 131807 4527 131835
rect 4561 131807 4589 131835
rect 4623 131807 4651 131835
rect 4437 131745 4465 131773
rect 4499 131745 4527 131773
rect 4561 131745 4589 131773
rect 4623 131745 4651 131773
rect 4437 122931 4465 122959
rect 4499 122931 4527 122959
rect 4561 122931 4589 122959
rect 4623 122931 4651 122959
rect 4437 122869 4465 122897
rect 4499 122869 4527 122897
rect 4561 122869 4589 122897
rect 4623 122869 4651 122897
rect 4437 122807 4465 122835
rect 4499 122807 4527 122835
rect 4561 122807 4589 122835
rect 4623 122807 4651 122835
rect 4437 122745 4465 122773
rect 4499 122745 4527 122773
rect 4561 122745 4589 122773
rect 4623 122745 4651 122773
rect 4437 113931 4465 113959
rect 4499 113931 4527 113959
rect 4561 113931 4589 113959
rect 4623 113931 4651 113959
rect 4437 113869 4465 113897
rect 4499 113869 4527 113897
rect 4561 113869 4589 113897
rect 4623 113869 4651 113897
rect 4437 113807 4465 113835
rect 4499 113807 4527 113835
rect 4561 113807 4589 113835
rect 4623 113807 4651 113835
rect 4437 113745 4465 113773
rect 4499 113745 4527 113773
rect 4561 113745 4589 113773
rect 4623 113745 4651 113773
rect 4437 104931 4465 104959
rect 4499 104931 4527 104959
rect 4561 104931 4589 104959
rect 4623 104931 4651 104959
rect 4437 104869 4465 104897
rect 4499 104869 4527 104897
rect 4561 104869 4589 104897
rect 4623 104869 4651 104897
rect 4437 104807 4465 104835
rect 4499 104807 4527 104835
rect 4561 104807 4589 104835
rect 4623 104807 4651 104835
rect 4437 104745 4465 104773
rect 4499 104745 4527 104773
rect 4561 104745 4589 104773
rect 4623 104745 4651 104773
rect 4437 95931 4465 95959
rect 4499 95931 4527 95959
rect 4561 95931 4589 95959
rect 4623 95931 4651 95959
rect 4437 95869 4465 95897
rect 4499 95869 4527 95897
rect 4561 95869 4589 95897
rect 4623 95869 4651 95897
rect 4437 95807 4465 95835
rect 4499 95807 4527 95835
rect 4561 95807 4589 95835
rect 4623 95807 4651 95835
rect 4437 95745 4465 95773
rect 4499 95745 4527 95773
rect 4561 95745 4589 95773
rect 4623 95745 4651 95773
rect 4437 86931 4465 86959
rect 4499 86931 4527 86959
rect 4561 86931 4589 86959
rect 4623 86931 4651 86959
rect 4437 86869 4465 86897
rect 4499 86869 4527 86897
rect 4561 86869 4589 86897
rect 4623 86869 4651 86897
rect 4437 86807 4465 86835
rect 4499 86807 4527 86835
rect 4561 86807 4589 86835
rect 4623 86807 4651 86835
rect 4437 86745 4465 86773
rect 4499 86745 4527 86773
rect 4561 86745 4589 86773
rect 4623 86745 4651 86773
rect 4437 77931 4465 77959
rect 4499 77931 4527 77959
rect 4561 77931 4589 77959
rect 4623 77931 4651 77959
rect 4437 77869 4465 77897
rect 4499 77869 4527 77897
rect 4561 77869 4589 77897
rect 4623 77869 4651 77897
rect 4437 77807 4465 77835
rect 4499 77807 4527 77835
rect 4561 77807 4589 77835
rect 4623 77807 4651 77835
rect 4437 77745 4465 77773
rect 4499 77745 4527 77773
rect 4561 77745 4589 77773
rect 4623 77745 4651 77773
rect 4437 68931 4465 68959
rect 4499 68931 4527 68959
rect 4561 68931 4589 68959
rect 4623 68931 4651 68959
rect 4437 68869 4465 68897
rect 4499 68869 4527 68897
rect 4561 68869 4589 68897
rect 4623 68869 4651 68897
rect 4437 68807 4465 68835
rect 4499 68807 4527 68835
rect 4561 68807 4589 68835
rect 4623 68807 4651 68835
rect 4437 68745 4465 68773
rect 4499 68745 4527 68773
rect 4561 68745 4589 68773
rect 4623 68745 4651 68773
rect 4437 59931 4465 59959
rect 4499 59931 4527 59959
rect 4561 59931 4589 59959
rect 4623 59931 4651 59959
rect 4437 59869 4465 59897
rect 4499 59869 4527 59897
rect 4561 59869 4589 59897
rect 4623 59869 4651 59897
rect 4437 59807 4465 59835
rect 4499 59807 4527 59835
rect 4561 59807 4589 59835
rect 4623 59807 4651 59835
rect 4437 59745 4465 59773
rect 4499 59745 4527 59773
rect 4561 59745 4589 59773
rect 4623 59745 4651 59773
rect 4437 50931 4465 50959
rect 4499 50931 4527 50959
rect 4561 50931 4589 50959
rect 4623 50931 4651 50959
rect 4437 50869 4465 50897
rect 4499 50869 4527 50897
rect 4561 50869 4589 50897
rect 4623 50869 4651 50897
rect 4437 50807 4465 50835
rect 4499 50807 4527 50835
rect 4561 50807 4589 50835
rect 4623 50807 4651 50835
rect 4437 50745 4465 50773
rect 4499 50745 4527 50773
rect 4561 50745 4589 50773
rect 4623 50745 4651 50773
rect 4437 41931 4465 41959
rect 4499 41931 4527 41959
rect 4561 41931 4589 41959
rect 4623 41931 4651 41959
rect 4437 41869 4465 41897
rect 4499 41869 4527 41897
rect 4561 41869 4589 41897
rect 4623 41869 4651 41897
rect 4437 41807 4465 41835
rect 4499 41807 4527 41835
rect 4561 41807 4589 41835
rect 4623 41807 4651 41835
rect 4437 41745 4465 41773
rect 4499 41745 4527 41773
rect 4561 41745 4589 41773
rect 4623 41745 4651 41773
rect 4437 32931 4465 32959
rect 4499 32931 4527 32959
rect 4561 32931 4589 32959
rect 4623 32931 4651 32959
rect 4437 32869 4465 32897
rect 4499 32869 4527 32897
rect 4561 32869 4589 32897
rect 4623 32869 4651 32897
rect 4437 32807 4465 32835
rect 4499 32807 4527 32835
rect 4561 32807 4589 32835
rect 4623 32807 4651 32835
rect 4437 32745 4465 32773
rect 4499 32745 4527 32773
rect 4561 32745 4589 32773
rect 4623 32745 4651 32773
rect 4437 23931 4465 23959
rect 4499 23931 4527 23959
rect 4561 23931 4589 23959
rect 4623 23931 4651 23959
rect 4437 23869 4465 23897
rect 4499 23869 4527 23897
rect 4561 23869 4589 23897
rect 4623 23869 4651 23897
rect 4437 23807 4465 23835
rect 4499 23807 4527 23835
rect 4561 23807 4589 23835
rect 4623 23807 4651 23835
rect 4437 23745 4465 23773
rect 4499 23745 4527 23773
rect 4561 23745 4589 23773
rect 4623 23745 4651 23773
rect 4437 14931 4465 14959
rect 4499 14931 4527 14959
rect 4561 14931 4589 14959
rect 4623 14931 4651 14959
rect 4437 14869 4465 14897
rect 4499 14869 4527 14897
rect 4561 14869 4589 14897
rect 4623 14869 4651 14897
rect 4437 14807 4465 14835
rect 4499 14807 4527 14835
rect 4561 14807 4589 14835
rect 4623 14807 4651 14835
rect 4437 14745 4465 14773
rect 4499 14745 4527 14773
rect 4561 14745 4589 14773
rect 4623 14745 4651 14773
rect 4437 5931 4465 5959
rect 4499 5931 4527 5959
rect 4561 5931 4589 5959
rect 4623 5931 4651 5959
rect 4437 5869 4465 5897
rect 4499 5869 4527 5897
rect 4561 5869 4589 5897
rect 4623 5869 4651 5897
rect 4437 5807 4465 5835
rect 4499 5807 4527 5835
rect 4561 5807 4589 5835
rect 4623 5807 4651 5835
rect 4437 5745 4465 5773
rect 4499 5745 4527 5773
rect 4561 5745 4589 5773
rect 4623 5745 4651 5773
rect 4437 396 4465 424
rect 4499 396 4527 424
rect 4561 396 4589 424
rect 4623 396 4651 424
rect 4437 334 4465 362
rect 4499 334 4527 362
rect 4561 334 4589 362
rect 4623 334 4651 362
rect 4437 272 4465 300
rect 4499 272 4527 300
rect 4561 272 4589 300
rect 4623 272 4651 300
rect 4437 210 4465 238
rect 4499 210 4527 238
rect 4561 210 4589 238
rect 4623 210 4651 238
rect 11577 299162 11605 299190
rect 11639 299162 11667 299190
rect 11701 299162 11729 299190
rect 11763 299162 11791 299190
rect 11577 299100 11605 299128
rect 11639 299100 11667 299128
rect 11701 299100 11729 299128
rect 11763 299100 11791 299128
rect 11577 299038 11605 299066
rect 11639 299038 11667 299066
rect 11701 299038 11729 299066
rect 11763 299038 11791 299066
rect 11577 298976 11605 299004
rect 11639 298976 11667 299004
rect 11701 298976 11729 299004
rect 11763 298976 11791 299004
rect 11577 290931 11605 290959
rect 11639 290931 11667 290959
rect 11701 290931 11729 290959
rect 11763 290931 11791 290959
rect 11577 290869 11605 290897
rect 11639 290869 11667 290897
rect 11701 290869 11729 290897
rect 11763 290869 11791 290897
rect 11577 290807 11605 290835
rect 11639 290807 11667 290835
rect 11701 290807 11729 290835
rect 11763 290807 11791 290835
rect 11577 290745 11605 290773
rect 11639 290745 11667 290773
rect 11701 290745 11729 290773
rect 11763 290745 11791 290773
rect 11577 281931 11605 281959
rect 11639 281931 11667 281959
rect 11701 281931 11729 281959
rect 11763 281931 11791 281959
rect 11577 281869 11605 281897
rect 11639 281869 11667 281897
rect 11701 281869 11729 281897
rect 11763 281869 11791 281897
rect 11577 281807 11605 281835
rect 11639 281807 11667 281835
rect 11701 281807 11729 281835
rect 11763 281807 11791 281835
rect 11577 281745 11605 281773
rect 11639 281745 11667 281773
rect 11701 281745 11729 281773
rect 11763 281745 11791 281773
rect 11577 272931 11605 272959
rect 11639 272931 11667 272959
rect 11701 272931 11729 272959
rect 11763 272931 11791 272959
rect 11577 272869 11605 272897
rect 11639 272869 11667 272897
rect 11701 272869 11729 272897
rect 11763 272869 11791 272897
rect 11577 272807 11605 272835
rect 11639 272807 11667 272835
rect 11701 272807 11729 272835
rect 11763 272807 11791 272835
rect 11577 272745 11605 272773
rect 11639 272745 11667 272773
rect 11701 272745 11729 272773
rect 11763 272745 11791 272773
rect 11577 263931 11605 263959
rect 11639 263931 11667 263959
rect 11701 263931 11729 263959
rect 11763 263931 11791 263959
rect 11577 263869 11605 263897
rect 11639 263869 11667 263897
rect 11701 263869 11729 263897
rect 11763 263869 11791 263897
rect 11577 263807 11605 263835
rect 11639 263807 11667 263835
rect 11701 263807 11729 263835
rect 11763 263807 11791 263835
rect 11577 263745 11605 263773
rect 11639 263745 11667 263773
rect 11701 263745 11729 263773
rect 11763 263745 11791 263773
rect 11577 254931 11605 254959
rect 11639 254931 11667 254959
rect 11701 254931 11729 254959
rect 11763 254931 11791 254959
rect 11577 254869 11605 254897
rect 11639 254869 11667 254897
rect 11701 254869 11729 254897
rect 11763 254869 11791 254897
rect 11577 254807 11605 254835
rect 11639 254807 11667 254835
rect 11701 254807 11729 254835
rect 11763 254807 11791 254835
rect 11577 254745 11605 254773
rect 11639 254745 11667 254773
rect 11701 254745 11729 254773
rect 11763 254745 11791 254773
rect 11577 245931 11605 245959
rect 11639 245931 11667 245959
rect 11701 245931 11729 245959
rect 11763 245931 11791 245959
rect 11577 245869 11605 245897
rect 11639 245869 11667 245897
rect 11701 245869 11729 245897
rect 11763 245869 11791 245897
rect 11577 245807 11605 245835
rect 11639 245807 11667 245835
rect 11701 245807 11729 245835
rect 11763 245807 11791 245835
rect 11577 245745 11605 245773
rect 11639 245745 11667 245773
rect 11701 245745 11729 245773
rect 11763 245745 11791 245773
rect 11577 236931 11605 236959
rect 11639 236931 11667 236959
rect 11701 236931 11729 236959
rect 11763 236931 11791 236959
rect 11577 236869 11605 236897
rect 11639 236869 11667 236897
rect 11701 236869 11729 236897
rect 11763 236869 11791 236897
rect 11577 236807 11605 236835
rect 11639 236807 11667 236835
rect 11701 236807 11729 236835
rect 11763 236807 11791 236835
rect 11577 236745 11605 236773
rect 11639 236745 11667 236773
rect 11701 236745 11729 236773
rect 11763 236745 11791 236773
rect 11577 227931 11605 227959
rect 11639 227931 11667 227959
rect 11701 227931 11729 227959
rect 11763 227931 11791 227959
rect 11577 227869 11605 227897
rect 11639 227869 11667 227897
rect 11701 227869 11729 227897
rect 11763 227869 11791 227897
rect 11577 227807 11605 227835
rect 11639 227807 11667 227835
rect 11701 227807 11729 227835
rect 11763 227807 11791 227835
rect 11577 227745 11605 227773
rect 11639 227745 11667 227773
rect 11701 227745 11729 227773
rect 11763 227745 11791 227773
rect 11577 218931 11605 218959
rect 11639 218931 11667 218959
rect 11701 218931 11729 218959
rect 11763 218931 11791 218959
rect 11577 218869 11605 218897
rect 11639 218869 11667 218897
rect 11701 218869 11729 218897
rect 11763 218869 11791 218897
rect 11577 218807 11605 218835
rect 11639 218807 11667 218835
rect 11701 218807 11729 218835
rect 11763 218807 11791 218835
rect 11577 218745 11605 218773
rect 11639 218745 11667 218773
rect 11701 218745 11729 218773
rect 11763 218745 11791 218773
rect 11577 209931 11605 209959
rect 11639 209931 11667 209959
rect 11701 209931 11729 209959
rect 11763 209931 11791 209959
rect 11577 209869 11605 209897
rect 11639 209869 11667 209897
rect 11701 209869 11729 209897
rect 11763 209869 11791 209897
rect 11577 209807 11605 209835
rect 11639 209807 11667 209835
rect 11701 209807 11729 209835
rect 11763 209807 11791 209835
rect 11577 209745 11605 209773
rect 11639 209745 11667 209773
rect 11701 209745 11729 209773
rect 11763 209745 11791 209773
rect 11577 200931 11605 200959
rect 11639 200931 11667 200959
rect 11701 200931 11729 200959
rect 11763 200931 11791 200959
rect 11577 200869 11605 200897
rect 11639 200869 11667 200897
rect 11701 200869 11729 200897
rect 11763 200869 11791 200897
rect 11577 200807 11605 200835
rect 11639 200807 11667 200835
rect 11701 200807 11729 200835
rect 11763 200807 11791 200835
rect 11577 200745 11605 200773
rect 11639 200745 11667 200773
rect 11701 200745 11729 200773
rect 11763 200745 11791 200773
rect 11577 191931 11605 191959
rect 11639 191931 11667 191959
rect 11701 191931 11729 191959
rect 11763 191931 11791 191959
rect 11577 191869 11605 191897
rect 11639 191869 11667 191897
rect 11701 191869 11729 191897
rect 11763 191869 11791 191897
rect 11577 191807 11605 191835
rect 11639 191807 11667 191835
rect 11701 191807 11729 191835
rect 11763 191807 11791 191835
rect 11577 191745 11605 191773
rect 11639 191745 11667 191773
rect 11701 191745 11729 191773
rect 11763 191745 11791 191773
rect 11577 182931 11605 182959
rect 11639 182931 11667 182959
rect 11701 182931 11729 182959
rect 11763 182931 11791 182959
rect 11577 182869 11605 182897
rect 11639 182869 11667 182897
rect 11701 182869 11729 182897
rect 11763 182869 11791 182897
rect 11577 182807 11605 182835
rect 11639 182807 11667 182835
rect 11701 182807 11729 182835
rect 11763 182807 11791 182835
rect 11577 182745 11605 182773
rect 11639 182745 11667 182773
rect 11701 182745 11729 182773
rect 11763 182745 11791 182773
rect 11577 173931 11605 173959
rect 11639 173931 11667 173959
rect 11701 173931 11729 173959
rect 11763 173931 11791 173959
rect 11577 173869 11605 173897
rect 11639 173869 11667 173897
rect 11701 173869 11729 173897
rect 11763 173869 11791 173897
rect 11577 173807 11605 173835
rect 11639 173807 11667 173835
rect 11701 173807 11729 173835
rect 11763 173807 11791 173835
rect 11577 173745 11605 173773
rect 11639 173745 11667 173773
rect 11701 173745 11729 173773
rect 11763 173745 11791 173773
rect 11577 164931 11605 164959
rect 11639 164931 11667 164959
rect 11701 164931 11729 164959
rect 11763 164931 11791 164959
rect 11577 164869 11605 164897
rect 11639 164869 11667 164897
rect 11701 164869 11729 164897
rect 11763 164869 11791 164897
rect 11577 164807 11605 164835
rect 11639 164807 11667 164835
rect 11701 164807 11729 164835
rect 11763 164807 11791 164835
rect 11577 164745 11605 164773
rect 11639 164745 11667 164773
rect 11701 164745 11729 164773
rect 11763 164745 11791 164773
rect 11577 155931 11605 155959
rect 11639 155931 11667 155959
rect 11701 155931 11729 155959
rect 11763 155931 11791 155959
rect 11577 155869 11605 155897
rect 11639 155869 11667 155897
rect 11701 155869 11729 155897
rect 11763 155869 11791 155897
rect 11577 155807 11605 155835
rect 11639 155807 11667 155835
rect 11701 155807 11729 155835
rect 11763 155807 11791 155835
rect 11577 155745 11605 155773
rect 11639 155745 11667 155773
rect 11701 155745 11729 155773
rect 11763 155745 11791 155773
rect 11577 146931 11605 146959
rect 11639 146931 11667 146959
rect 11701 146931 11729 146959
rect 11763 146931 11791 146959
rect 11577 146869 11605 146897
rect 11639 146869 11667 146897
rect 11701 146869 11729 146897
rect 11763 146869 11791 146897
rect 11577 146807 11605 146835
rect 11639 146807 11667 146835
rect 11701 146807 11729 146835
rect 11763 146807 11791 146835
rect 11577 146745 11605 146773
rect 11639 146745 11667 146773
rect 11701 146745 11729 146773
rect 11763 146745 11791 146773
rect 11577 137931 11605 137959
rect 11639 137931 11667 137959
rect 11701 137931 11729 137959
rect 11763 137931 11791 137959
rect 11577 137869 11605 137897
rect 11639 137869 11667 137897
rect 11701 137869 11729 137897
rect 11763 137869 11791 137897
rect 11577 137807 11605 137835
rect 11639 137807 11667 137835
rect 11701 137807 11729 137835
rect 11763 137807 11791 137835
rect 11577 137745 11605 137773
rect 11639 137745 11667 137773
rect 11701 137745 11729 137773
rect 11763 137745 11791 137773
rect 11577 128931 11605 128959
rect 11639 128931 11667 128959
rect 11701 128931 11729 128959
rect 11763 128931 11791 128959
rect 11577 128869 11605 128897
rect 11639 128869 11667 128897
rect 11701 128869 11729 128897
rect 11763 128869 11791 128897
rect 11577 128807 11605 128835
rect 11639 128807 11667 128835
rect 11701 128807 11729 128835
rect 11763 128807 11791 128835
rect 11577 128745 11605 128773
rect 11639 128745 11667 128773
rect 11701 128745 11729 128773
rect 11763 128745 11791 128773
rect 11577 119931 11605 119959
rect 11639 119931 11667 119959
rect 11701 119931 11729 119959
rect 11763 119931 11791 119959
rect 11577 119869 11605 119897
rect 11639 119869 11667 119897
rect 11701 119869 11729 119897
rect 11763 119869 11791 119897
rect 11577 119807 11605 119835
rect 11639 119807 11667 119835
rect 11701 119807 11729 119835
rect 11763 119807 11791 119835
rect 11577 119745 11605 119773
rect 11639 119745 11667 119773
rect 11701 119745 11729 119773
rect 11763 119745 11791 119773
rect 11577 110931 11605 110959
rect 11639 110931 11667 110959
rect 11701 110931 11729 110959
rect 11763 110931 11791 110959
rect 11577 110869 11605 110897
rect 11639 110869 11667 110897
rect 11701 110869 11729 110897
rect 11763 110869 11791 110897
rect 11577 110807 11605 110835
rect 11639 110807 11667 110835
rect 11701 110807 11729 110835
rect 11763 110807 11791 110835
rect 11577 110745 11605 110773
rect 11639 110745 11667 110773
rect 11701 110745 11729 110773
rect 11763 110745 11791 110773
rect 11577 101931 11605 101959
rect 11639 101931 11667 101959
rect 11701 101931 11729 101959
rect 11763 101931 11791 101959
rect 11577 101869 11605 101897
rect 11639 101869 11667 101897
rect 11701 101869 11729 101897
rect 11763 101869 11791 101897
rect 11577 101807 11605 101835
rect 11639 101807 11667 101835
rect 11701 101807 11729 101835
rect 11763 101807 11791 101835
rect 11577 101745 11605 101773
rect 11639 101745 11667 101773
rect 11701 101745 11729 101773
rect 11763 101745 11791 101773
rect 11577 92931 11605 92959
rect 11639 92931 11667 92959
rect 11701 92931 11729 92959
rect 11763 92931 11791 92959
rect 11577 92869 11605 92897
rect 11639 92869 11667 92897
rect 11701 92869 11729 92897
rect 11763 92869 11791 92897
rect 11577 92807 11605 92835
rect 11639 92807 11667 92835
rect 11701 92807 11729 92835
rect 11763 92807 11791 92835
rect 11577 92745 11605 92773
rect 11639 92745 11667 92773
rect 11701 92745 11729 92773
rect 11763 92745 11791 92773
rect 11577 83931 11605 83959
rect 11639 83931 11667 83959
rect 11701 83931 11729 83959
rect 11763 83931 11791 83959
rect 11577 83869 11605 83897
rect 11639 83869 11667 83897
rect 11701 83869 11729 83897
rect 11763 83869 11791 83897
rect 11577 83807 11605 83835
rect 11639 83807 11667 83835
rect 11701 83807 11729 83835
rect 11763 83807 11791 83835
rect 11577 83745 11605 83773
rect 11639 83745 11667 83773
rect 11701 83745 11729 83773
rect 11763 83745 11791 83773
rect 11577 74931 11605 74959
rect 11639 74931 11667 74959
rect 11701 74931 11729 74959
rect 11763 74931 11791 74959
rect 11577 74869 11605 74897
rect 11639 74869 11667 74897
rect 11701 74869 11729 74897
rect 11763 74869 11791 74897
rect 11577 74807 11605 74835
rect 11639 74807 11667 74835
rect 11701 74807 11729 74835
rect 11763 74807 11791 74835
rect 11577 74745 11605 74773
rect 11639 74745 11667 74773
rect 11701 74745 11729 74773
rect 11763 74745 11791 74773
rect 11577 65931 11605 65959
rect 11639 65931 11667 65959
rect 11701 65931 11729 65959
rect 11763 65931 11791 65959
rect 11577 65869 11605 65897
rect 11639 65869 11667 65897
rect 11701 65869 11729 65897
rect 11763 65869 11791 65897
rect 11577 65807 11605 65835
rect 11639 65807 11667 65835
rect 11701 65807 11729 65835
rect 11763 65807 11791 65835
rect 11577 65745 11605 65773
rect 11639 65745 11667 65773
rect 11701 65745 11729 65773
rect 11763 65745 11791 65773
rect 11577 56931 11605 56959
rect 11639 56931 11667 56959
rect 11701 56931 11729 56959
rect 11763 56931 11791 56959
rect 11577 56869 11605 56897
rect 11639 56869 11667 56897
rect 11701 56869 11729 56897
rect 11763 56869 11791 56897
rect 11577 56807 11605 56835
rect 11639 56807 11667 56835
rect 11701 56807 11729 56835
rect 11763 56807 11791 56835
rect 11577 56745 11605 56773
rect 11639 56745 11667 56773
rect 11701 56745 11729 56773
rect 11763 56745 11791 56773
rect 11577 47931 11605 47959
rect 11639 47931 11667 47959
rect 11701 47931 11729 47959
rect 11763 47931 11791 47959
rect 11577 47869 11605 47897
rect 11639 47869 11667 47897
rect 11701 47869 11729 47897
rect 11763 47869 11791 47897
rect 11577 47807 11605 47835
rect 11639 47807 11667 47835
rect 11701 47807 11729 47835
rect 11763 47807 11791 47835
rect 11577 47745 11605 47773
rect 11639 47745 11667 47773
rect 11701 47745 11729 47773
rect 11763 47745 11791 47773
rect 11577 38931 11605 38959
rect 11639 38931 11667 38959
rect 11701 38931 11729 38959
rect 11763 38931 11791 38959
rect 11577 38869 11605 38897
rect 11639 38869 11667 38897
rect 11701 38869 11729 38897
rect 11763 38869 11791 38897
rect 11577 38807 11605 38835
rect 11639 38807 11667 38835
rect 11701 38807 11729 38835
rect 11763 38807 11791 38835
rect 11577 38745 11605 38773
rect 11639 38745 11667 38773
rect 11701 38745 11729 38773
rect 11763 38745 11791 38773
rect 11577 29931 11605 29959
rect 11639 29931 11667 29959
rect 11701 29931 11729 29959
rect 11763 29931 11791 29959
rect 11577 29869 11605 29897
rect 11639 29869 11667 29897
rect 11701 29869 11729 29897
rect 11763 29869 11791 29897
rect 11577 29807 11605 29835
rect 11639 29807 11667 29835
rect 11701 29807 11729 29835
rect 11763 29807 11791 29835
rect 11577 29745 11605 29773
rect 11639 29745 11667 29773
rect 11701 29745 11729 29773
rect 11763 29745 11791 29773
rect 11577 20931 11605 20959
rect 11639 20931 11667 20959
rect 11701 20931 11729 20959
rect 11763 20931 11791 20959
rect 11577 20869 11605 20897
rect 11639 20869 11667 20897
rect 11701 20869 11729 20897
rect 11763 20869 11791 20897
rect 11577 20807 11605 20835
rect 11639 20807 11667 20835
rect 11701 20807 11729 20835
rect 11763 20807 11791 20835
rect 11577 20745 11605 20773
rect 11639 20745 11667 20773
rect 11701 20745 11729 20773
rect 11763 20745 11791 20773
rect 11577 11931 11605 11959
rect 11639 11931 11667 11959
rect 11701 11931 11729 11959
rect 11763 11931 11791 11959
rect 11577 11869 11605 11897
rect 11639 11869 11667 11897
rect 11701 11869 11729 11897
rect 11763 11869 11791 11897
rect 11577 11807 11605 11835
rect 11639 11807 11667 11835
rect 11701 11807 11729 11835
rect 11763 11807 11791 11835
rect 11577 11745 11605 11773
rect 11639 11745 11667 11773
rect 11701 11745 11729 11773
rect 11763 11745 11791 11773
rect 11577 2931 11605 2959
rect 11639 2931 11667 2959
rect 11701 2931 11729 2959
rect 11763 2931 11791 2959
rect 11577 2869 11605 2897
rect 11639 2869 11667 2897
rect 11701 2869 11729 2897
rect 11763 2869 11791 2897
rect 11577 2807 11605 2835
rect 11639 2807 11667 2835
rect 11701 2807 11729 2835
rect 11763 2807 11791 2835
rect 11577 2745 11605 2773
rect 11639 2745 11667 2773
rect 11701 2745 11729 2773
rect 11763 2745 11791 2773
rect 11577 876 11605 904
rect 11639 876 11667 904
rect 11701 876 11729 904
rect 11763 876 11791 904
rect 11577 814 11605 842
rect 11639 814 11667 842
rect 11701 814 11729 842
rect 11763 814 11791 842
rect 11577 752 11605 780
rect 11639 752 11667 780
rect 11701 752 11729 780
rect 11763 752 11791 780
rect 11577 690 11605 718
rect 11639 690 11667 718
rect 11701 690 11729 718
rect 11763 690 11791 718
rect 13437 299642 13465 299670
rect 13499 299642 13527 299670
rect 13561 299642 13589 299670
rect 13623 299642 13651 299670
rect 13437 299580 13465 299608
rect 13499 299580 13527 299608
rect 13561 299580 13589 299608
rect 13623 299580 13651 299608
rect 13437 299518 13465 299546
rect 13499 299518 13527 299546
rect 13561 299518 13589 299546
rect 13623 299518 13651 299546
rect 13437 299456 13465 299484
rect 13499 299456 13527 299484
rect 13561 299456 13589 299484
rect 13623 299456 13651 299484
rect 13437 293931 13465 293959
rect 13499 293931 13527 293959
rect 13561 293931 13589 293959
rect 13623 293931 13651 293959
rect 13437 293869 13465 293897
rect 13499 293869 13527 293897
rect 13561 293869 13589 293897
rect 13623 293869 13651 293897
rect 13437 293807 13465 293835
rect 13499 293807 13527 293835
rect 13561 293807 13589 293835
rect 13623 293807 13651 293835
rect 13437 293745 13465 293773
rect 13499 293745 13527 293773
rect 13561 293745 13589 293773
rect 13623 293745 13651 293773
rect 13437 284931 13465 284959
rect 13499 284931 13527 284959
rect 13561 284931 13589 284959
rect 13623 284931 13651 284959
rect 13437 284869 13465 284897
rect 13499 284869 13527 284897
rect 13561 284869 13589 284897
rect 13623 284869 13651 284897
rect 13437 284807 13465 284835
rect 13499 284807 13527 284835
rect 13561 284807 13589 284835
rect 13623 284807 13651 284835
rect 13437 284745 13465 284773
rect 13499 284745 13527 284773
rect 13561 284745 13589 284773
rect 13623 284745 13651 284773
rect 13437 275931 13465 275959
rect 13499 275931 13527 275959
rect 13561 275931 13589 275959
rect 13623 275931 13651 275959
rect 13437 275869 13465 275897
rect 13499 275869 13527 275897
rect 13561 275869 13589 275897
rect 13623 275869 13651 275897
rect 13437 275807 13465 275835
rect 13499 275807 13527 275835
rect 13561 275807 13589 275835
rect 13623 275807 13651 275835
rect 13437 275745 13465 275773
rect 13499 275745 13527 275773
rect 13561 275745 13589 275773
rect 13623 275745 13651 275773
rect 13437 266931 13465 266959
rect 13499 266931 13527 266959
rect 13561 266931 13589 266959
rect 13623 266931 13651 266959
rect 13437 266869 13465 266897
rect 13499 266869 13527 266897
rect 13561 266869 13589 266897
rect 13623 266869 13651 266897
rect 13437 266807 13465 266835
rect 13499 266807 13527 266835
rect 13561 266807 13589 266835
rect 13623 266807 13651 266835
rect 13437 266745 13465 266773
rect 13499 266745 13527 266773
rect 13561 266745 13589 266773
rect 13623 266745 13651 266773
rect 13437 257931 13465 257959
rect 13499 257931 13527 257959
rect 13561 257931 13589 257959
rect 13623 257931 13651 257959
rect 13437 257869 13465 257897
rect 13499 257869 13527 257897
rect 13561 257869 13589 257897
rect 13623 257869 13651 257897
rect 13437 257807 13465 257835
rect 13499 257807 13527 257835
rect 13561 257807 13589 257835
rect 13623 257807 13651 257835
rect 13437 257745 13465 257773
rect 13499 257745 13527 257773
rect 13561 257745 13589 257773
rect 13623 257745 13651 257773
rect 20577 299162 20605 299190
rect 20639 299162 20667 299190
rect 20701 299162 20729 299190
rect 20763 299162 20791 299190
rect 20577 299100 20605 299128
rect 20639 299100 20667 299128
rect 20701 299100 20729 299128
rect 20763 299100 20791 299128
rect 20577 299038 20605 299066
rect 20639 299038 20667 299066
rect 20701 299038 20729 299066
rect 20763 299038 20791 299066
rect 20577 298976 20605 299004
rect 20639 298976 20667 299004
rect 20701 298976 20729 299004
rect 20763 298976 20791 299004
rect 20577 290931 20605 290959
rect 20639 290931 20667 290959
rect 20701 290931 20729 290959
rect 20763 290931 20791 290959
rect 20577 290869 20605 290897
rect 20639 290869 20667 290897
rect 20701 290869 20729 290897
rect 20763 290869 20791 290897
rect 20577 290807 20605 290835
rect 20639 290807 20667 290835
rect 20701 290807 20729 290835
rect 20763 290807 20791 290835
rect 20577 290745 20605 290773
rect 20639 290745 20667 290773
rect 20701 290745 20729 290773
rect 20763 290745 20791 290773
rect 20577 281931 20605 281959
rect 20639 281931 20667 281959
rect 20701 281931 20729 281959
rect 20763 281931 20791 281959
rect 20577 281869 20605 281897
rect 20639 281869 20667 281897
rect 20701 281869 20729 281897
rect 20763 281869 20791 281897
rect 20577 281807 20605 281835
rect 20639 281807 20667 281835
rect 20701 281807 20729 281835
rect 20763 281807 20791 281835
rect 20577 281745 20605 281773
rect 20639 281745 20667 281773
rect 20701 281745 20729 281773
rect 20763 281745 20791 281773
rect 20577 272931 20605 272959
rect 20639 272931 20667 272959
rect 20701 272931 20729 272959
rect 20763 272931 20791 272959
rect 20577 272869 20605 272897
rect 20639 272869 20667 272897
rect 20701 272869 20729 272897
rect 20763 272869 20791 272897
rect 20577 272807 20605 272835
rect 20639 272807 20667 272835
rect 20701 272807 20729 272835
rect 20763 272807 20791 272835
rect 20577 272745 20605 272773
rect 20639 272745 20667 272773
rect 20701 272745 20729 272773
rect 20763 272745 20791 272773
rect 20577 263931 20605 263959
rect 20639 263931 20667 263959
rect 20701 263931 20729 263959
rect 20763 263931 20791 263959
rect 20577 263869 20605 263897
rect 20639 263869 20667 263897
rect 20701 263869 20729 263897
rect 20763 263869 20791 263897
rect 20577 263807 20605 263835
rect 20639 263807 20667 263835
rect 20701 263807 20729 263835
rect 20763 263807 20791 263835
rect 20577 263745 20605 263773
rect 20639 263745 20667 263773
rect 20701 263745 20729 263773
rect 20763 263745 20791 263773
rect 20577 254931 20605 254959
rect 20639 254931 20667 254959
rect 20701 254931 20729 254959
rect 20763 254931 20791 254959
rect 20577 254869 20605 254897
rect 20639 254869 20667 254897
rect 20701 254869 20729 254897
rect 20763 254869 20791 254897
rect 20577 254807 20605 254835
rect 20639 254807 20667 254835
rect 20701 254807 20729 254835
rect 20763 254807 20791 254835
rect 20577 254745 20605 254773
rect 20639 254745 20667 254773
rect 20701 254745 20729 254773
rect 20763 254745 20791 254773
rect 13437 248931 13465 248959
rect 13499 248931 13527 248959
rect 13561 248931 13589 248959
rect 13623 248931 13651 248959
rect 13437 248869 13465 248897
rect 13499 248869 13527 248897
rect 13561 248869 13589 248897
rect 13623 248869 13651 248897
rect 13437 248807 13465 248835
rect 13499 248807 13527 248835
rect 13561 248807 13589 248835
rect 13623 248807 13651 248835
rect 13437 248745 13465 248773
rect 13499 248745 13527 248773
rect 13561 248745 13589 248773
rect 13623 248745 13651 248773
rect 17259 245931 17287 245959
rect 17321 245931 17349 245959
rect 17259 245869 17287 245897
rect 17321 245869 17349 245897
rect 17259 245807 17287 245835
rect 17321 245807 17349 245835
rect 17259 245745 17287 245773
rect 17321 245745 17349 245773
rect 20577 245931 20605 245959
rect 20639 245931 20667 245959
rect 20701 245931 20729 245959
rect 20763 245931 20791 245959
rect 20577 245869 20605 245897
rect 20639 245869 20667 245897
rect 20701 245869 20729 245897
rect 20763 245869 20791 245897
rect 20577 245807 20605 245835
rect 20639 245807 20667 245835
rect 20701 245807 20729 245835
rect 20763 245807 20791 245835
rect 20577 245745 20605 245773
rect 20639 245745 20667 245773
rect 20701 245745 20729 245773
rect 20763 245745 20791 245773
rect 13437 239931 13465 239959
rect 13499 239931 13527 239959
rect 13561 239931 13589 239959
rect 13623 239931 13651 239959
rect 13437 239869 13465 239897
rect 13499 239869 13527 239897
rect 13561 239869 13589 239897
rect 13623 239869 13651 239897
rect 13437 239807 13465 239835
rect 13499 239807 13527 239835
rect 13561 239807 13589 239835
rect 13623 239807 13651 239835
rect 13437 239745 13465 239773
rect 13499 239745 13527 239773
rect 13561 239745 13589 239773
rect 13623 239745 13651 239773
rect 17259 236931 17287 236959
rect 17321 236931 17349 236959
rect 17259 236869 17287 236897
rect 17321 236869 17349 236897
rect 17259 236807 17287 236835
rect 17321 236807 17349 236835
rect 17259 236745 17287 236773
rect 17321 236745 17349 236773
rect 20577 236931 20605 236959
rect 20639 236931 20667 236959
rect 20701 236931 20729 236959
rect 20763 236931 20791 236959
rect 20577 236869 20605 236897
rect 20639 236869 20667 236897
rect 20701 236869 20729 236897
rect 20763 236869 20791 236897
rect 20577 236807 20605 236835
rect 20639 236807 20667 236835
rect 20701 236807 20729 236835
rect 20763 236807 20791 236835
rect 20577 236745 20605 236773
rect 20639 236745 20667 236773
rect 20701 236745 20729 236773
rect 20763 236745 20791 236773
rect 13437 230931 13465 230959
rect 13499 230931 13527 230959
rect 13561 230931 13589 230959
rect 13623 230931 13651 230959
rect 13437 230869 13465 230897
rect 13499 230869 13527 230897
rect 13561 230869 13589 230897
rect 13623 230869 13651 230897
rect 13437 230807 13465 230835
rect 13499 230807 13527 230835
rect 13561 230807 13589 230835
rect 13623 230807 13651 230835
rect 13437 230745 13465 230773
rect 13499 230745 13527 230773
rect 13561 230745 13589 230773
rect 13623 230745 13651 230773
rect 17259 227931 17287 227959
rect 17321 227931 17349 227959
rect 17259 227869 17287 227897
rect 17321 227869 17349 227897
rect 17259 227807 17287 227835
rect 17321 227807 17349 227835
rect 17259 227745 17287 227773
rect 17321 227745 17349 227773
rect 20577 227931 20605 227959
rect 20639 227931 20667 227959
rect 20701 227931 20729 227959
rect 20763 227931 20791 227959
rect 20577 227869 20605 227897
rect 20639 227869 20667 227897
rect 20701 227869 20729 227897
rect 20763 227869 20791 227897
rect 20577 227807 20605 227835
rect 20639 227807 20667 227835
rect 20701 227807 20729 227835
rect 20763 227807 20791 227835
rect 20577 227745 20605 227773
rect 20639 227745 20667 227773
rect 20701 227745 20729 227773
rect 20763 227745 20791 227773
rect 13437 221931 13465 221959
rect 13499 221931 13527 221959
rect 13561 221931 13589 221959
rect 13623 221931 13651 221959
rect 13437 221869 13465 221897
rect 13499 221869 13527 221897
rect 13561 221869 13589 221897
rect 13623 221869 13651 221897
rect 13437 221807 13465 221835
rect 13499 221807 13527 221835
rect 13561 221807 13589 221835
rect 13623 221807 13651 221835
rect 13437 221745 13465 221773
rect 13499 221745 13527 221773
rect 13561 221745 13589 221773
rect 13623 221745 13651 221773
rect 17259 218931 17287 218959
rect 17321 218931 17349 218959
rect 17259 218869 17287 218897
rect 17321 218869 17349 218897
rect 17259 218807 17287 218835
rect 17321 218807 17349 218835
rect 17259 218745 17287 218773
rect 17321 218745 17349 218773
rect 20577 218931 20605 218959
rect 20639 218931 20667 218959
rect 20701 218931 20729 218959
rect 20763 218931 20791 218959
rect 20577 218869 20605 218897
rect 20639 218869 20667 218897
rect 20701 218869 20729 218897
rect 20763 218869 20791 218897
rect 20577 218807 20605 218835
rect 20639 218807 20667 218835
rect 20701 218807 20729 218835
rect 20763 218807 20791 218835
rect 20577 218745 20605 218773
rect 20639 218745 20667 218773
rect 20701 218745 20729 218773
rect 20763 218745 20791 218773
rect 13437 212931 13465 212959
rect 13499 212931 13527 212959
rect 13561 212931 13589 212959
rect 13623 212931 13651 212959
rect 13437 212869 13465 212897
rect 13499 212869 13527 212897
rect 13561 212869 13589 212897
rect 13623 212869 13651 212897
rect 13437 212807 13465 212835
rect 13499 212807 13527 212835
rect 13561 212807 13589 212835
rect 13623 212807 13651 212835
rect 13437 212745 13465 212773
rect 13499 212745 13527 212773
rect 13561 212745 13589 212773
rect 13623 212745 13651 212773
rect 17259 209931 17287 209959
rect 17321 209931 17349 209959
rect 17259 209869 17287 209897
rect 17321 209869 17349 209897
rect 17259 209807 17287 209835
rect 17321 209807 17349 209835
rect 17259 209745 17287 209773
rect 17321 209745 17349 209773
rect 20577 209931 20605 209959
rect 20639 209931 20667 209959
rect 20701 209931 20729 209959
rect 20763 209931 20791 209959
rect 20577 209869 20605 209897
rect 20639 209869 20667 209897
rect 20701 209869 20729 209897
rect 20763 209869 20791 209897
rect 20577 209807 20605 209835
rect 20639 209807 20667 209835
rect 20701 209807 20729 209835
rect 20763 209807 20791 209835
rect 20577 209745 20605 209773
rect 20639 209745 20667 209773
rect 20701 209745 20729 209773
rect 20763 209745 20791 209773
rect 13437 203931 13465 203959
rect 13499 203931 13527 203959
rect 13561 203931 13589 203959
rect 13623 203931 13651 203959
rect 13437 203869 13465 203897
rect 13499 203869 13527 203897
rect 13561 203869 13589 203897
rect 13623 203869 13651 203897
rect 13437 203807 13465 203835
rect 13499 203807 13527 203835
rect 13561 203807 13589 203835
rect 13623 203807 13651 203835
rect 13437 203745 13465 203773
rect 13499 203745 13527 203773
rect 13561 203745 13589 203773
rect 13623 203745 13651 203773
rect 17259 200931 17287 200959
rect 17321 200931 17349 200959
rect 17259 200869 17287 200897
rect 17321 200869 17349 200897
rect 17259 200807 17287 200835
rect 17321 200807 17349 200835
rect 17259 200745 17287 200773
rect 17321 200745 17349 200773
rect 20577 200931 20605 200959
rect 20639 200931 20667 200959
rect 20701 200931 20729 200959
rect 20763 200931 20791 200959
rect 20577 200869 20605 200897
rect 20639 200869 20667 200897
rect 20701 200869 20729 200897
rect 20763 200869 20791 200897
rect 20577 200807 20605 200835
rect 20639 200807 20667 200835
rect 20701 200807 20729 200835
rect 20763 200807 20791 200835
rect 20577 200745 20605 200773
rect 20639 200745 20667 200773
rect 20701 200745 20729 200773
rect 20763 200745 20791 200773
rect 13437 194931 13465 194959
rect 13499 194931 13527 194959
rect 13561 194931 13589 194959
rect 13623 194931 13651 194959
rect 13437 194869 13465 194897
rect 13499 194869 13527 194897
rect 13561 194869 13589 194897
rect 13623 194869 13651 194897
rect 13437 194807 13465 194835
rect 13499 194807 13527 194835
rect 13561 194807 13589 194835
rect 13623 194807 13651 194835
rect 13437 194745 13465 194773
rect 13499 194745 13527 194773
rect 13561 194745 13589 194773
rect 13623 194745 13651 194773
rect 17259 191931 17287 191959
rect 17321 191931 17349 191959
rect 17259 191869 17287 191897
rect 17321 191869 17349 191897
rect 17259 191807 17287 191835
rect 17321 191807 17349 191835
rect 17259 191745 17287 191773
rect 17321 191745 17349 191773
rect 20577 191931 20605 191959
rect 20639 191931 20667 191959
rect 20701 191931 20729 191959
rect 20763 191931 20791 191959
rect 20577 191869 20605 191897
rect 20639 191869 20667 191897
rect 20701 191869 20729 191897
rect 20763 191869 20791 191897
rect 20577 191807 20605 191835
rect 20639 191807 20667 191835
rect 20701 191807 20729 191835
rect 20763 191807 20791 191835
rect 20577 191745 20605 191773
rect 20639 191745 20667 191773
rect 20701 191745 20729 191773
rect 20763 191745 20791 191773
rect 13437 185931 13465 185959
rect 13499 185931 13527 185959
rect 13561 185931 13589 185959
rect 13623 185931 13651 185959
rect 13437 185869 13465 185897
rect 13499 185869 13527 185897
rect 13561 185869 13589 185897
rect 13623 185869 13651 185897
rect 13437 185807 13465 185835
rect 13499 185807 13527 185835
rect 13561 185807 13589 185835
rect 13623 185807 13651 185835
rect 13437 185745 13465 185773
rect 13499 185745 13527 185773
rect 13561 185745 13589 185773
rect 13623 185745 13651 185773
rect 17259 182931 17287 182959
rect 17321 182931 17349 182959
rect 17259 182869 17287 182897
rect 17321 182869 17349 182897
rect 17259 182807 17287 182835
rect 17321 182807 17349 182835
rect 17259 182745 17287 182773
rect 17321 182745 17349 182773
rect 20577 182931 20605 182959
rect 20639 182931 20667 182959
rect 20701 182931 20729 182959
rect 20763 182931 20791 182959
rect 20577 182869 20605 182897
rect 20639 182869 20667 182897
rect 20701 182869 20729 182897
rect 20763 182869 20791 182897
rect 20577 182807 20605 182835
rect 20639 182807 20667 182835
rect 20701 182807 20729 182835
rect 20763 182807 20791 182835
rect 20577 182745 20605 182773
rect 20639 182745 20667 182773
rect 20701 182745 20729 182773
rect 20763 182745 20791 182773
rect 13437 176931 13465 176959
rect 13499 176931 13527 176959
rect 13561 176931 13589 176959
rect 13623 176931 13651 176959
rect 13437 176869 13465 176897
rect 13499 176869 13527 176897
rect 13561 176869 13589 176897
rect 13623 176869 13651 176897
rect 13437 176807 13465 176835
rect 13499 176807 13527 176835
rect 13561 176807 13589 176835
rect 13623 176807 13651 176835
rect 13437 176745 13465 176773
rect 13499 176745 13527 176773
rect 13561 176745 13589 176773
rect 13623 176745 13651 176773
rect 17259 173931 17287 173959
rect 17321 173931 17349 173959
rect 17259 173869 17287 173897
rect 17321 173869 17349 173897
rect 17259 173807 17287 173835
rect 17321 173807 17349 173835
rect 17259 173745 17287 173773
rect 17321 173745 17349 173773
rect 20577 173931 20605 173959
rect 20639 173931 20667 173959
rect 20701 173931 20729 173959
rect 20763 173931 20791 173959
rect 20577 173869 20605 173897
rect 20639 173869 20667 173897
rect 20701 173869 20729 173897
rect 20763 173869 20791 173897
rect 20577 173807 20605 173835
rect 20639 173807 20667 173835
rect 20701 173807 20729 173835
rect 20763 173807 20791 173835
rect 20577 173745 20605 173773
rect 20639 173745 20667 173773
rect 20701 173745 20729 173773
rect 20763 173745 20791 173773
rect 13437 167931 13465 167959
rect 13499 167931 13527 167959
rect 13561 167931 13589 167959
rect 13623 167931 13651 167959
rect 13437 167869 13465 167897
rect 13499 167869 13527 167897
rect 13561 167869 13589 167897
rect 13623 167869 13651 167897
rect 13437 167807 13465 167835
rect 13499 167807 13527 167835
rect 13561 167807 13589 167835
rect 13623 167807 13651 167835
rect 13437 167745 13465 167773
rect 13499 167745 13527 167773
rect 13561 167745 13589 167773
rect 13623 167745 13651 167773
rect 17259 164931 17287 164959
rect 17321 164931 17349 164959
rect 17259 164869 17287 164897
rect 17321 164869 17349 164897
rect 17259 164807 17287 164835
rect 17321 164807 17349 164835
rect 17259 164745 17287 164773
rect 17321 164745 17349 164773
rect 20577 164931 20605 164959
rect 20639 164931 20667 164959
rect 20701 164931 20729 164959
rect 20763 164931 20791 164959
rect 20577 164869 20605 164897
rect 20639 164869 20667 164897
rect 20701 164869 20729 164897
rect 20763 164869 20791 164897
rect 20577 164807 20605 164835
rect 20639 164807 20667 164835
rect 20701 164807 20729 164835
rect 20763 164807 20791 164835
rect 20577 164745 20605 164773
rect 20639 164745 20667 164773
rect 20701 164745 20729 164773
rect 20763 164745 20791 164773
rect 13437 158931 13465 158959
rect 13499 158931 13527 158959
rect 13561 158931 13589 158959
rect 13623 158931 13651 158959
rect 13437 158869 13465 158897
rect 13499 158869 13527 158897
rect 13561 158869 13589 158897
rect 13623 158869 13651 158897
rect 13437 158807 13465 158835
rect 13499 158807 13527 158835
rect 13561 158807 13589 158835
rect 13623 158807 13651 158835
rect 13437 158745 13465 158773
rect 13499 158745 13527 158773
rect 13561 158745 13589 158773
rect 13623 158745 13651 158773
rect 17259 155931 17287 155959
rect 17321 155931 17349 155959
rect 17259 155869 17287 155897
rect 17321 155869 17349 155897
rect 17259 155807 17287 155835
rect 17321 155807 17349 155835
rect 17259 155745 17287 155773
rect 17321 155745 17349 155773
rect 20577 155931 20605 155959
rect 20639 155931 20667 155959
rect 20701 155931 20729 155959
rect 20763 155931 20791 155959
rect 20577 155869 20605 155897
rect 20639 155869 20667 155897
rect 20701 155869 20729 155897
rect 20763 155869 20791 155897
rect 20577 155807 20605 155835
rect 20639 155807 20667 155835
rect 20701 155807 20729 155835
rect 20763 155807 20791 155835
rect 20577 155745 20605 155773
rect 20639 155745 20667 155773
rect 20701 155745 20729 155773
rect 20763 155745 20791 155773
rect 13437 149931 13465 149959
rect 13499 149931 13527 149959
rect 13561 149931 13589 149959
rect 13623 149931 13651 149959
rect 13437 149869 13465 149897
rect 13499 149869 13527 149897
rect 13561 149869 13589 149897
rect 13623 149869 13651 149897
rect 13437 149807 13465 149835
rect 13499 149807 13527 149835
rect 13561 149807 13589 149835
rect 13623 149807 13651 149835
rect 13437 149745 13465 149773
rect 13499 149745 13527 149773
rect 13561 149745 13589 149773
rect 13623 149745 13651 149773
rect 17259 146931 17287 146959
rect 17321 146931 17349 146959
rect 17259 146869 17287 146897
rect 17321 146869 17349 146897
rect 17259 146807 17287 146835
rect 17321 146807 17349 146835
rect 17259 146745 17287 146773
rect 17321 146745 17349 146773
rect 20577 146931 20605 146959
rect 20639 146931 20667 146959
rect 20701 146931 20729 146959
rect 20763 146931 20791 146959
rect 20577 146869 20605 146897
rect 20639 146869 20667 146897
rect 20701 146869 20729 146897
rect 20763 146869 20791 146897
rect 20577 146807 20605 146835
rect 20639 146807 20667 146835
rect 20701 146807 20729 146835
rect 20763 146807 20791 146835
rect 20577 146745 20605 146773
rect 20639 146745 20667 146773
rect 20701 146745 20729 146773
rect 20763 146745 20791 146773
rect 13437 140931 13465 140959
rect 13499 140931 13527 140959
rect 13561 140931 13589 140959
rect 13623 140931 13651 140959
rect 13437 140869 13465 140897
rect 13499 140869 13527 140897
rect 13561 140869 13589 140897
rect 13623 140869 13651 140897
rect 13437 140807 13465 140835
rect 13499 140807 13527 140835
rect 13561 140807 13589 140835
rect 13623 140807 13651 140835
rect 13437 140745 13465 140773
rect 13499 140745 13527 140773
rect 13561 140745 13589 140773
rect 13623 140745 13651 140773
rect 17259 137931 17287 137959
rect 17321 137931 17349 137959
rect 17259 137869 17287 137897
rect 17321 137869 17349 137897
rect 17259 137807 17287 137835
rect 17321 137807 17349 137835
rect 17259 137745 17287 137773
rect 17321 137745 17349 137773
rect 20577 137931 20605 137959
rect 20639 137931 20667 137959
rect 20701 137931 20729 137959
rect 20763 137931 20791 137959
rect 20577 137869 20605 137897
rect 20639 137869 20667 137897
rect 20701 137869 20729 137897
rect 20763 137869 20791 137897
rect 20577 137807 20605 137835
rect 20639 137807 20667 137835
rect 20701 137807 20729 137835
rect 20763 137807 20791 137835
rect 20577 137745 20605 137773
rect 20639 137745 20667 137773
rect 20701 137745 20729 137773
rect 20763 137745 20791 137773
rect 13437 131931 13465 131959
rect 13499 131931 13527 131959
rect 13561 131931 13589 131959
rect 13623 131931 13651 131959
rect 13437 131869 13465 131897
rect 13499 131869 13527 131897
rect 13561 131869 13589 131897
rect 13623 131869 13651 131897
rect 13437 131807 13465 131835
rect 13499 131807 13527 131835
rect 13561 131807 13589 131835
rect 13623 131807 13651 131835
rect 13437 131745 13465 131773
rect 13499 131745 13527 131773
rect 13561 131745 13589 131773
rect 13623 131745 13651 131773
rect 17259 128931 17287 128959
rect 17321 128931 17349 128959
rect 17259 128869 17287 128897
rect 17321 128869 17349 128897
rect 17259 128807 17287 128835
rect 17321 128807 17349 128835
rect 17259 128745 17287 128773
rect 17321 128745 17349 128773
rect 20577 128931 20605 128959
rect 20639 128931 20667 128959
rect 20701 128931 20729 128959
rect 20763 128931 20791 128959
rect 20577 128869 20605 128897
rect 20639 128869 20667 128897
rect 20701 128869 20729 128897
rect 20763 128869 20791 128897
rect 20577 128807 20605 128835
rect 20639 128807 20667 128835
rect 20701 128807 20729 128835
rect 20763 128807 20791 128835
rect 20577 128745 20605 128773
rect 20639 128745 20667 128773
rect 20701 128745 20729 128773
rect 20763 128745 20791 128773
rect 13437 122931 13465 122959
rect 13499 122931 13527 122959
rect 13561 122931 13589 122959
rect 13623 122931 13651 122959
rect 13437 122869 13465 122897
rect 13499 122869 13527 122897
rect 13561 122869 13589 122897
rect 13623 122869 13651 122897
rect 13437 122807 13465 122835
rect 13499 122807 13527 122835
rect 13561 122807 13589 122835
rect 13623 122807 13651 122835
rect 13437 122745 13465 122773
rect 13499 122745 13527 122773
rect 13561 122745 13589 122773
rect 13623 122745 13651 122773
rect 17259 119931 17287 119959
rect 17321 119931 17349 119959
rect 17259 119869 17287 119897
rect 17321 119869 17349 119897
rect 17259 119807 17287 119835
rect 17321 119807 17349 119835
rect 17259 119745 17287 119773
rect 17321 119745 17349 119773
rect 20577 119931 20605 119959
rect 20639 119931 20667 119959
rect 20701 119931 20729 119959
rect 20763 119931 20791 119959
rect 20577 119869 20605 119897
rect 20639 119869 20667 119897
rect 20701 119869 20729 119897
rect 20763 119869 20791 119897
rect 20577 119807 20605 119835
rect 20639 119807 20667 119835
rect 20701 119807 20729 119835
rect 20763 119807 20791 119835
rect 20577 119745 20605 119773
rect 20639 119745 20667 119773
rect 20701 119745 20729 119773
rect 20763 119745 20791 119773
rect 13437 113931 13465 113959
rect 13499 113931 13527 113959
rect 13561 113931 13589 113959
rect 13623 113931 13651 113959
rect 13437 113869 13465 113897
rect 13499 113869 13527 113897
rect 13561 113869 13589 113897
rect 13623 113869 13651 113897
rect 13437 113807 13465 113835
rect 13499 113807 13527 113835
rect 13561 113807 13589 113835
rect 13623 113807 13651 113835
rect 13437 113745 13465 113773
rect 13499 113745 13527 113773
rect 13561 113745 13589 113773
rect 13623 113745 13651 113773
rect 17259 110931 17287 110959
rect 17321 110931 17349 110959
rect 17259 110869 17287 110897
rect 17321 110869 17349 110897
rect 17259 110807 17287 110835
rect 17321 110807 17349 110835
rect 17259 110745 17287 110773
rect 17321 110745 17349 110773
rect 20577 110931 20605 110959
rect 20639 110931 20667 110959
rect 20701 110931 20729 110959
rect 20763 110931 20791 110959
rect 20577 110869 20605 110897
rect 20639 110869 20667 110897
rect 20701 110869 20729 110897
rect 20763 110869 20791 110897
rect 20577 110807 20605 110835
rect 20639 110807 20667 110835
rect 20701 110807 20729 110835
rect 20763 110807 20791 110835
rect 20577 110745 20605 110773
rect 20639 110745 20667 110773
rect 20701 110745 20729 110773
rect 20763 110745 20791 110773
rect 13437 104931 13465 104959
rect 13499 104931 13527 104959
rect 13561 104931 13589 104959
rect 13623 104931 13651 104959
rect 13437 104869 13465 104897
rect 13499 104869 13527 104897
rect 13561 104869 13589 104897
rect 13623 104869 13651 104897
rect 13437 104807 13465 104835
rect 13499 104807 13527 104835
rect 13561 104807 13589 104835
rect 13623 104807 13651 104835
rect 13437 104745 13465 104773
rect 13499 104745 13527 104773
rect 13561 104745 13589 104773
rect 13623 104745 13651 104773
rect 17259 101931 17287 101959
rect 17321 101931 17349 101959
rect 17259 101869 17287 101897
rect 17321 101869 17349 101897
rect 17259 101807 17287 101835
rect 17321 101807 17349 101835
rect 17259 101745 17287 101773
rect 17321 101745 17349 101773
rect 20577 101931 20605 101959
rect 20639 101931 20667 101959
rect 20701 101931 20729 101959
rect 20763 101931 20791 101959
rect 20577 101869 20605 101897
rect 20639 101869 20667 101897
rect 20701 101869 20729 101897
rect 20763 101869 20791 101897
rect 20577 101807 20605 101835
rect 20639 101807 20667 101835
rect 20701 101807 20729 101835
rect 20763 101807 20791 101835
rect 20577 101745 20605 101773
rect 20639 101745 20667 101773
rect 20701 101745 20729 101773
rect 20763 101745 20791 101773
rect 13437 95931 13465 95959
rect 13499 95931 13527 95959
rect 13561 95931 13589 95959
rect 13623 95931 13651 95959
rect 13437 95869 13465 95897
rect 13499 95869 13527 95897
rect 13561 95869 13589 95897
rect 13623 95869 13651 95897
rect 13437 95807 13465 95835
rect 13499 95807 13527 95835
rect 13561 95807 13589 95835
rect 13623 95807 13651 95835
rect 13437 95745 13465 95773
rect 13499 95745 13527 95773
rect 13561 95745 13589 95773
rect 13623 95745 13651 95773
rect 17259 92931 17287 92959
rect 17321 92931 17349 92959
rect 17259 92869 17287 92897
rect 17321 92869 17349 92897
rect 17259 92807 17287 92835
rect 17321 92807 17349 92835
rect 17259 92745 17287 92773
rect 17321 92745 17349 92773
rect 20577 92931 20605 92959
rect 20639 92931 20667 92959
rect 20701 92931 20729 92959
rect 20763 92931 20791 92959
rect 20577 92869 20605 92897
rect 20639 92869 20667 92897
rect 20701 92869 20729 92897
rect 20763 92869 20791 92897
rect 20577 92807 20605 92835
rect 20639 92807 20667 92835
rect 20701 92807 20729 92835
rect 20763 92807 20791 92835
rect 20577 92745 20605 92773
rect 20639 92745 20667 92773
rect 20701 92745 20729 92773
rect 20763 92745 20791 92773
rect 13437 86931 13465 86959
rect 13499 86931 13527 86959
rect 13561 86931 13589 86959
rect 13623 86931 13651 86959
rect 13437 86869 13465 86897
rect 13499 86869 13527 86897
rect 13561 86869 13589 86897
rect 13623 86869 13651 86897
rect 13437 86807 13465 86835
rect 13499 86807 13527 86835
rect 13561 86807 13589 86835
rect 13623 86807 13651 86835
rect 13437 86745 13465 86773
rect 13499 86745 13527 86773
rect 13561 86745 13589 86773
rect 13623 86745 13651 86773
rect 17259 83931 17287 83959
rect 17321 83931 17349 83959
rect 17259 83869 17287 83897
rect 17321 83869 17349 83897
rect 17259 83807 17287 83835
rect 17321 83807 17349 83835
rect 17259 83745 17287 83773
rect 17321 83745 17349 83773
rect 20577 83931 20605 83959
rect 20639 83931 20667 83959
rect 20701 83931 20729 83959
rect 20763 83931 20791 83959
rect 20577 83869 20605 83897
rect 20639 83869 20667 83897
rect 20701 83869 20729 83897
rect 20763 83869 20791 83897
rect 20577 83807 20605 83835
rect 20639 83807 20667 83835
rect 20701 83807 20729 83835
rect 20763 83807 20791 83835
rect 20577 83745 20605 83773
rect 20639 83745 20667 83773
rect 20701 83745 20729 83773
rect 20763 83745 20791 83773
rect 13437 77931 13465 77959
rect 13499 77931 13527 77959
rect 13561 77931 13589 77959
rect 13623 77931 13651 77959
rect 13437 77869 13465 77897
rect 13499 77869 13527 77897
rect 13561 77869 13589 77897
rect 13623 77869 13651 77897
rect 13437 77807 13465 77835
rect 13499 77807 13527 77835
rect 13561 77807 13589 77835
rect 13623 77807 13651 77835
rect 13437 77745 13465 77773
rect 13499 77745 13527 77773
rect 13561 77745 13589 77773
rect 13623 77745 13651 77773
rect 17259 74931 17287 74959
rect 17321 74931 17349 74959
rect 17259 74869 17287 74897
rect 17321 74869 17349 74897
rect 17259 74807 17287 74835
rect 17321 74807 17349 74835
rect 17259 74745 17287 74773
rect 17321 74745 17349 74773
rect 20577 74931 20605 74959
rect 20639 74931 20667 74959
rect 20701 74931 20729 74959
rect 20763 74931 20791 74959
rect 20577 74869 20605 74897
rect 20639 74869 20667 74897
rect 20701 74869 20729 74897
rect 20763 74869 20791 74897
rect 20577 74807 20605 74835
rect 20639 74807 20667 74835
rect 20701 74807 20729 74835
rect 20763 74807 20791 74835
rect 20577 74745 20605 74773
rect 20639 74745 20667 74773
rect 20701 74745 20729 74773
rect 20763 74745 20791 74773
rect 13437 68931 13465 68959
rect 13499 68931 13527 68959
rect 13561 68931 13589 68959
rect 13623 68931 13651 68959
rect 13437 68869 13465 68897
rect 13499 68869 13527 68897
rect 13561 68869 13589 68897
rect 13623 68869 13651 68897
rect 13437 68807 13465 68835
rect 13499 68807 13527 68835
rect 13561 68807 13589 68835
rect 13623 68807 13651 68835
rect 13437 68745 13465 68773
rect 13499 68745 13527 68773
rect 13561 68745 13589 68773
rect 13623 68745 13651 68773
rect 17259 65931 17287 65959
rect 17321 65931 17349 65959
rect 17259 65869 17287 65897
rect 17321 65869 17349 65897
rect 17259 65807 17287 65835
rect 17321 65807 17349 65835
rect 17259 65745 17287 65773
rect 17321 65745 17349 65773
rect 20577 65931 20605 65959
rect 20639 65931 20667 65959
rect 20701 65931 20729 65959
rect 20763 65931 20791 65959
rect 20577 65869 20605 65897
rect 20639 65869 20667 65897
rect 20701 65869 20729 65897
rect 20763 65869 20791 65897
rect 20577 65807 20605 65835
rect 20639 65807 20667 65835
rect 20701 65807 20729 65835
rect 20763 65807 20791 65835
rect 20577 65745 20605 65773
rect 20639 65745 20667 65773
rect 20701 65745 20729 65773
rect 20763 65745 20791 65773
rect 13437 59931 13465 59959
rect 13499 59931 13527 59959
rect 13561 59931 13589 59959
rect 13623 59931 13651 59959
rect 13437 59869 13465 59897
rect 13499 59869 13527 59897
rect 13561 59869 13589 59897
rect 13623 59869 13651 59897
rect 13437 59807 13465 59835
rect 13499 59807 13527 59835
rect 13561 59807 13589 59835
rect 13623 59807 13651 59835
rect 13437 59745 13465 59773
rect 13499 59745 13527 59773
rect 13561 59745 13589 59773
rect 13623 59745 13651 59773
rect 17259 56931 17287 56959
rect 17321 56931 17349 56959
rect 17259 56869 17287 56897
rect 17321 56869 17349 56897
rect 17259 56807 17287 56835
rect 17321 56807 17349 56835
rect 17259 56745 17287 56773
rect 17321 56745 17349 56773
rect 20577 56931 20605 56959
rect 20639 56931 20667 56959
rect 20701 56931 20729 56959
rect 20763 56931 20791 56959
rect 20577 56869 20605 56897
rect 20639 56869 20667 56897
rect 20701 56869 20729 56897
rect 20763 56869 20791 56897
rect 20577 56807 20605 56835
rect 20639 56807 20667 56835
rect 20701 56807 20729 56835
rect 20763 56807 20791 56835
rect 20577 56745 20605 56773
rect 20639 56745 20667 56773
rect 20701 56745 20729 56773
rect 20763 56745 20791 56773
rect 13437 50931 13465 50959
rect 13499 50931 13527 50959
rect 13561 50931 13589 50959
rect 13623 50931 13651 50959
rect 13437 50869 13465 50897
rect 13499 50869 13527 50897
rect 13561 50869 13589 50897
rect 13623 50869 13651 50897
rect 13437 50807 13465 50835
rect 13499 50807 13527 50835
rect 13561 50807 13589 50835
rect 13623 50807 13651 50835
rect 13437 50745 13465 50773
rect 13499 50745 13527 50773
rect 13561 50745 13589 50773
rect 13623 50745 13651 50773
rect 17259 47931 17287 47959
rect 17321 47931 17349 47959
rect 17259 47869 17287 47897
rect 17321 47869 17349 47897
rect 17259 47807 17287 47835
rect 17321 47807 17349 47835
rect 17259 47745 17287 47773
rect 17321 47745 17349 47773
rect 20577 47931 20605 47959
rect 20639 47931 20667 47959
rect 20701 47931 20729 47959
rect 20763 47931 20791 47959
rect 20577 47869 20605 47897
rect 20639 47869 20667 47897
rect 20701 47869 20729 47897
rect 20763 47869 20791 47897
rect 20577 47807 20605 47835
rect 20639 47807 20667 47835
rect 20701 47807 20729 47835
rect 20763 47807 20791 47835
rect 20577 47745 20605 47773
rect 20639 47745 20667 47773
rect 20701 47745 20729 47773
rect 20763 47745 20791 47773
rect 13437 41931 13465 41959
rect 13499 41931 13527 41959
rect 13561 41931 13589 41959
rect 13623 41931 13651 41959
rect 13437 41869 13465 41897
rect 13499 41869 13527 41897
rect 13561 41869 13589 41897
rect 13623 41869 13651 41897
rect 13437 41807 13465 41835
rect 13499 41807 13527 41835
rect 13561 41807 13589 41835
rect 13623 41807 13651 41835
rect 13437 41745 13465 41773
rect 13499 41745 13527 41773
rect 13561 41745 13589 41773
rect 13623 41745 13651 41773
rect 17259 38931 17287 38959
rect 17321 38931 17349 38959
rect 17259 38869 17287 38897
rect 17321 38869 17349 38897
rect 17259 38807 17287 38835
rect 17321 38807 17349 38835
rect 17259 38745 17287 38773
rect 17321 38745 17349 38773
rect 20577 38931 20605 38959
rect 20639 38931 20667 38959
rect 20701 38931 20729 38959
rect 20763 38931 20791 38959
rect 20577 38869 20605 38897
rect 20639 38869 20667 38897
rect 20701 38869 20729 38897
rect 20763 38869 20791 38897
rect 20577 38807 20605 38835
rect 20639 38807 20667 38835
rect 20701 38807 20729 38835
rect 20763 38807 20791 38835
rect 20577 38745 20605 38773
rect 20639 38745 20667 38773
rect 20701 38745 20729 38773
rect 20763 38745 20791 38773
rect 13437 32931 13465 32959
rect 13499 32931 13527 32959
rect 13561 32931 13589 32959
rect 13623 32931 13651 32959
rect 13437 32869 13465 32897
rect 13499 32869 13527 32897
rect 13561 32869 13589 32897
rect 13623 32869 13651 32897
rect 13437 32807 13465 32835
rect 13499 32807 13527 32835
rect 13561 32807 13589 32835
rect 13623 32807 13651 32835
rect 13437 32745 13465 32773
rect 13499 32745 13527 32773
rect 13561 32745 13589 32773
rect 13623 32745 13651 32773
rect 17259 29931 17287 29959
rect 17321 29931 17349 29959
rect 17259 29869 17287 29897
rect 17321 29869 17349 29897
rect 17259 29807 17287 29835
rect 17321 29807 17349 29835
rect 17259 29745 17287 29773
rect 17321 29745 17349 29773
rect 20577 29931 20605 29959
rect 20639 29931 20667 29959
rect 20701 29931 20729 29959
rect 20763 29931 20791 29959
rect 20577 29869 20605 29897
rect 20639 29869 20667 29897
rect 20701 29869 20729 29897
rect 20763 29869 20791 29897
rect 20577 29807 20605 29835
rect 20639 29807 20667 29835
rect 20701 29807 20729 29835
rect 20763 29807 20791 29835
rect 20577 29745 20605 29773
rect 20639 29745 20667 29773
rect 20701 29745 20729 29773
rect 20763 29745 20791 29773
rect 13437 23931 13465 23959
rect 13499 23931 13527 23959
rect 13561 23931 13589 23959
rect 13623 23931 13651 23959
rect 13437 23869 13465 23897
rect 13499 23869 13527 23897
rect 13561 23869 13589 23897
rect 13623 23869 13651 23897
rect 13437 23807 13465 23835
rect 13499 23807 13527 23835
rect 13561 23807 13589 23835
rect 13623 23807 13651 23835
rect 13437 23745 13465 23773
rect 13499 23745 13527 23773
rect 13561 23745 13589 23773
rect 13623 23745 13651 23773
rect 17259 20931 17287 20959
rect 17321 20931 17349 20959
rect 17259 20869 17287 20897
rect 17321 20869 17349 20897
rect 17259 20807 17287 20835
rect 17321 20807 17349 20835
rect 17259 20745 17287 20773
rect 17321 20745 17349 20773
rect 20577 20931 20605 20959
rect 20639 20931 20667 20959
rect 20701 20931 20729 20959
rect 20763 20931 20791 20959
rect 20577 20869 20605 20897
rect 20639 20869 20667 20897
rect 20701 20869 20729 20897
rect 20763 20869 20791 20897
rect 20577 20807 20605 20835
rect 20639 20807 20667 20835
rect 20701 20807 20729 20835
rect 20763 20807 20791 20835
rect 20577 20745 20605 20773
rect 20639 20745 20667 20773
rect 20701 20745 20729 20773
rect 20763 20745 20791 20773
rect 13437 14931 13465 14959
rect 13499 14931 13527 14959
rect 13561 14931 13589 14959
rect 13623 14931 13651 14959
rect 13437 14869 13465 14897
rect 13499 14869 13527 14897
rect 13561 14869 13589 14897
rect 13623 14869 13651 14897
rect 13437 14807 13465 14835
rect 13499 14807 13527 14835
rect 13561 14807 13589 14835
rect 13623 14807 13651 14835
rect 13437 14745 13465 14773
rect 13499 14745 13527 14773
rect 13561 14745 13589 14773
rect 13623 14745 13651 14773
rect 13437 5931 13465 5959
rect 13499 5931 13527 5959
rect 13561 5931 13589 5959
rect 13623 5931 13651 5959
rect 13437 5869 13465 5897
rect 13499 5869 13527 5897
rect 13561 5869 13589 5897
rect 13623 5869 13651 5897
rect 13437 5807 13465 5835
rect 13499 5807 13527 5835
rect 13561 5807 13589 5835
rect 13623 5807 13651 5835
rect 13437 5745 13465 5773
rect 13499 5745 13527 5773
rect 13561 5745 13589 5773
rect 13623 5745 13651 5773
rect 13437 396 13465 424
rect 13499 396 13527 424
rect 13561 396 13589 424
rect 13623 396 13651 424
rect 13437 334 13465 362
rect 13499 334 13527 362
rect 13561 334 13589 362
rect 13623 334 13651 362
rect 13437 272 13465 300
rect 13499 272 13527 300
rect 13561 272 13589 300
rect 13623 272 13651 300
rect 13437 210 13465 238
rect 13499 210 13527 238
rect 13561 210 13589 238
rect 13623 210 13651 238
rect 20577 11931 20605 11959
rect 20639 11931 20667 11959
rect 20701 11931 20729 11959
rect 20763 11931 20791 11959
rect 20577 11869 20605 11897
rect 20639 11869 20667 11897
rect 20701 11869 20729 11897
rect 20763 11869 20791 11897
rect 20577 11807 20605 11835
rect 20639 11807 20667 11835
rect 20701 11807 20729 11835
rect 20763 11807 20791 11835
rect 20577 11745 20605 11773
rect 20639 11745 20667 11773
rect 20701 11745 20729 11773
rect 20763 11745 20791 11773
rect 20577 2931 20605 2959
rect 20639 2931 20667 2959
rect 20701 2931 20729 2959
rect 20763 2931 20791 2959
rect 20577 2869 20605 2897
rect 20639 2869 20667 2897
rect 20701 2869 20729 2897
rect 20763 2869 20791 2897
rect 20577 2807 20605 2835
rect 20639 2807 20667 2835
rect 20701 2807 20729 2835
rect 20763 2807 20791 2835
rect 20577 2745 20605 2773
rect 20639 2745 20667 2773
rect 20701 2745 20729 2773
rect 20763 2745 20791 2773
rect 20577 876 20605 904
rect 20639 876 20667 904
rect 20701 876 20729 904
rect 20763 876 20791 904
rect 20577 814 20605 842
rect 20639 814 20667 842
rect 20701 814 20729 842
rect 20763 814 20791 842
rect 20577 752 20605 780
rect 20639 752 20667 780
rect 20701 752 20729 780
rect 20763 752 20791 780
rect 20577 690 20605 718
rect 20639 690 20667 718
rect 20701 690 20729 718
rect 20763 690 20791 718
rect 22437 299642 22465 299670
rect 22499 299642 22527 299670
rect 22561 299642 22589 299670
rect 22623 299642 22651 299670
rect 22437 299580 22465 299608
rect 22499 299580 22527 299608
rect 22561 299580 22589 299608
rect 22623 299580 22651 299608
rect 22437 299518 22465 299546
rect 22499 299518 22527 299546
rect 22561 299518 22589 299546
rect 22623 299518 22651 299546
rect 22437 299456 22465 299484
rect 22499 299456 22527 299484
rect 22561 299456 22589 299484
rect 22623 299456 22651 299484
rect 22437 293931 22465 293959
rect 22499 293931 22527 293959
rect 22561 293931 22589 293959
rect 22623 293931 22651 293959
rect 22437 293869 22465 293897
rect 22499 293869 22527 293897
rect 22561 293869 22589 293897
rect 22623 293869 22651 293897
rect 22437 293807 22465 293835
rect 22499 293807 22527 293835
rect 22561 293807 22589 293835
rect 22623 293807 22651 293835
rect 22437 293745 22465 293773
rect 22499 293745 22527 293773
rect 22561 293745 22589 293773
rect 22623 293745 22651 293773
rect 22437 284931 22465 284959
rect 22499 284931 22527 284959
rect 22561 284931 22589 284959
rect 22623 284931 22651 284959
rect 22437 284869 22465 284897
rect 22499 284869 22527 284897
rect 22561 284869 22589 284897
rect 22623 284869 22651 284897
rect 22437 284807 22465 284835
rect 22499 284807 22527 284835
rect 22561 284807 22589 284835
rect 22623 284807 22651 284835
rect 22437 284745 22465 284773
rect 22499 284745 22527 284773
rect 22561 284745 22589 284773
rect 22623 284745 22651 284773
rect 22437 275931 22465 275959
rect 22499 275931 22527 275959
rect 22561 275931 22589 275959
rect 22623 275931 22651 275959
rect 22437 275869 22465 275897
rect 22499 275869 22527 275897
rect 22561 275869 22589 275897
rect 22623 275869 22651 275897
rect 22437 275807 22465 275835
rect 22499 275807 22527 275835
rect 22561 275807 22589 275835
rect 22623 275807 22651 275835
rect 22437 275745 22465 275773
rect 22499 275745 22527 275773
rect 22561 275745 22589 275773
rect 22623 275745 22651 275773
rect 22437 266931 22465 266959
rect 22499 266931 22527 266959
rect 22561 266931 22589 266959
rect 22623 266931 22651 266959
rect 22437 266869 22465 266897
rect 22499 266869 22527 266897
rect 22561 266869 22589 266897
rect 22623 266869 22651 266897
rect 22437 266807 22465 266835
rect 22499 266807 22527 266835
rect 22561 266807 22589 266835
rect 22623 266807 22651 266835
rect 22437 266745 22465 266773
rect 22499 266745 22527 266773
rect 22561 266745 22589 266773
rect 22623 266745 22651 266773
rect 22437 257931 22465 257959
rect 22499 257931 22527 257959
rect 22561 257931 22589 257959
rect 22623 257931 22651 257959
rect 22437 257869 22465 257897
rect 22499 257869 22527 257897
rect 22561 257869 22589 257897
rect 22623 257869 22651 257897
rect 22437 257807 22465 257835
rect 22499 257807 22527 257835
rect 22561 257807 22589 257835
rect 22623 257807 22651 257835
rect 22437 257745 22465 257773
rect 22499 257745 22527 257773
rect 22561 257745 22589 257773
rect 22623 257745 22651 257773
rect 29577 299162 29605 299190
rect 29639 299162 29667 299190
rect 29701 299162 29729 299190
rect 29763 299162 29791 299190
rect 29577 299100 29605 299128
rect 29639 299100 29667 299128
rect 29701 299100 29729 299128
rect 29763 299100 29791 299128
rect 29577 299038 29605 299066
rect 29639 299038 29667 299066
rect 29701 299038 29729 299066
rect 29763 299038 29791 299066
rect 29577 298976 29605 299004
rect 29639 298976 29667 299004
rect 29701 298976 29729 299004
rect 29763 298976 29791 299004
rect 29577 290931 29605 290959
rect 29639 290931 29667 290959
rect 29701 290931 29729 290959
rect 29763 290931 29791 290959
rect 29577 290869 29605 290897
rect 29639 290869 29667 290897
rect 29701 290869 29729 290897
rect 29763 290869 29791 290897
rect 29577 290807 29605 290835
rect 29639 290807 29667 290835
rect 29701 290807 29729 290835
rect 29763 290807 29791 290835
rect 29577 290745 29605 290773
rect 29639 290745 29667 290773
rect 29701 290745 29729 290773
rect 29763 290745 29791 290773
rect 29577 281931 29605 281959
rect 29639 281931 29667 281959
rect 29701 281931 29729 281959
rect 29763 281931 29791 281959
rect 29577 281869 29605 281897
rect 29639 281869 29667 281897
rect 29701 281869 29729 281897
rect 29763 281869 29791 281897
rect 29577 281807 29605 281835
rect 29639 281807 29667 281835
rect 29701 281807 29729 281835
rect 29763 281807 29791 281835
rect 29577 281745 29605 281773
rect 29639 281745 29667 281773
rect 29701 281745 29729 281773
rect 29763 281745 29791 281773
rect 29577 272931 29605 272959
rect 29639 272931 29667 272959
rect 29701 272931 29729 272959
rect 29763 272931 29791 272959
rect 29577 272869 29605 272897
rect 29639 272869 29667 272897
rect 29701 272869 29729 272897
rect 29763 272869 29791 272897
rect 29577 272807 29605 272835
rect 29639 272807 29667 272835
rect 29701 272807 29729 272835
rect 29763 272807 29791 272835
rect 29577 272745 29605 272773
rect 29639 272745 29667 272773
rect 29701 272745 29729 272773
rect 29763 272745 29791 272773
rect 29577 263931 29605 263959
rect 29639 263931 29667 263959
rect 29701 263931 29729 263959
rect 29763 263931 29791 263959
rect 29577 263869 29605 263897
rect 29639 263869 29667 263897
rect 29701 263869 29729 263897
rect 29763 263869 29791 263897
rect 29577 263807 29605 263835
rect 29639 263807 29667 263835
rect 29701 263807 29729 263835
rect 29763 263807 29791 263835
rect 29577 263745 29605 263773
rect 29639 263745 29667 263773
rect 29701 263745 29729 263773
rect 29763 263745 29791 263773
rect 29577 254931 29605 254959
rect 29639 254931 29667 254959
rect 29701 254931 29729 254959
rect 29763 254931 29791 254959
rect 29577 254869 29605 254897
rect 29639 254869 29667 254897
rect 29701 254869 29729 254897
rect 29763 254869 29791 254897
rect 29577 254807 29605 254835
rect 29639 254807 29667 254835
rect 29701 254807 29729 254835
rect 29763 254807 29791 254835
rect 29577 254745 29605 254773
rect 29639 254745 29667 254773
rect 29701 254745 29729 254773
rect 29763 254745 29791 254773
rect 22437 248931 22465 248959
rect 22499 248931 22527 248959
rect 22561 248931 22589 248959
rect 22623 248931 22651 248959
rect 22437 248869 22465 248897
rect 22499 248869 22527 248897
rect 22561 248869 22589 248897
rect 22623 248869 22651 248897
rect 22437 248807 22465 248835
rect 22499 248807 22527 248835
rect 22561 248807 22589 248835
rect 22623 248807 22651 248835
rect 22437 248745 22465 248773
rect 22499 248745 22527 248773
rect 22561 248745 22589 248773
rect 22623 248745 22651 248773
rect 24939 248931 24967 248959
rect 25001 248931 25029 248959
rect 24939 248869 24967 248897
rect 25001 248869 25029 248897
rect 24939 248807 24967 248835
rect 25001 248807 25029 248835
rect 24939 248745 24967 248773
rect 25001 248745 25029 248773
rect 29577 245931 29605 245959
rect 29639 245931 29667 245959
rect 29701 245931 29729 245959
rect 29763 245931 29791 245959
rect 29577 245869 29605 245897
rect 29639 245869 29667 245897
rect 29701 245869 29729 245897
rect 29763 245869 29791 245897
rect 29577 245807 29605 245835
rect 29639 245807 29667 245835
rect 29701 245807 29729 245835
rect 29763 245807 29791 245835
rect 29577 245745 29605 245773
rect 29639 245745 29667 245773
rect 29701 245745 29729 245773
rect 29763 245745 29791 245773
rect 22437 239931 22465 239959
rect 22499 239931 22527 239959
rect 22561 239931 22589 239959
rect 22623 239931 22651 239959
rect 22437 239869 22465 239897
rect 22499 239869 22527 239897
rect 22561 239869 22589 239897
rect 22623 239869 22651 239897
rect 22437 239807 22465 239835
rect 22499 239807 22527 239835
rect 22561 239807 22589 239835
rect 22623 239807 22651 239835
rect 22437 239745 22465 239773
rect 22499 239745 22527 239773
rect 22561 239745 22589 239773
rect 22623 239745 22651 239773
rect 24939 239931 24967 239959
rect 25001 239931 25029 239959
rect 24939 239869 24967 239897
rect 25001 239869 25029 239897
rect 24939 239807 24967 239835
rect 25001 239807 25029 239835
rect 24939 239745 24967 239773
rect 25001 239745 25029 239773
rect 29577 236931 29605 236959
rect 29639 236931 29667 236959
rect 29701 236931 29729 236959
rect 29763 236931 29791 236959
rect 29577 236869 29605 236897
rect 29639 236869 29667 236897
rect 29701 236869 29729 236897
rect 29763 236869 29791 236897
rect 29577 236807 29605 236835
rect 29639 236807 29667 236835
rect 29701 236807 29729 236835
rect 29763 236807 29791 236835
rect 29577 236745 29605 236773
rect 29639 236745 29667 236773
rect 29701 236745 29729 236773
rect 29763 236745 29791 236773
rect 22437 230931 22465 230959
rect 22499 230931 22527 230959
rect 22561 230931 22589 230959
rect 22623 230931 22651 230959
rect 22437 230869 22465 230897
rect 22499 230869 22527 230897
rect 22561 230869 22589 230897
rect 22623 230869 22651 230897
rect 22437 230807 22465 230835
rect 22499 230807 22527 230835
rect 22561 230807 22589 230835
rect 22623 230807 22651 230835
rect 22437 230745 22465 230773
rect 22499 230745 22527 230773
rect 22561 230745 22589 230773
rect 22623 230745 22651 230773
rect 24939 230931 24967 230959
rect 25001 230931 25029 230959
rect 24939 230869 24967 230897
rect 25001 230869 25029 230897
rect 24939 230807 24967 230835
rect 25001 230807 25029 230835
rect 24939 230745 24967 230773
rect 25001 230745 25029 230773
rect 29577 227931 29605 227959
rect 29639 227931 29667 227959
rect 29701 227931 29729 227959
rect 29763 227931 29791 227959
rect 29577 227869 29605 227897
rect 29639 227869 29667 227897
rect 29701 227869 29729 227897
rect 29763 227869 29791 227897
rect 29577 227807 29605 227835
rect 29639 227807 29667 227835
rect 29701 227807 29729 227835
rect 29763 227807 29791 227835
rect 29577 227745 29605 227773
rect 29639 227745 29667 227773
rect 29701 227745 29729 227773
rect 29763 227745 29791 227773
rect 22437 221931 22465 221959
rect 22499 221931 22527 221959
rect 22561 221931 22589 221959
rect 22623 221931 22651 221959
rect 22437 221869 22465 221897
rect 22499 221869 22527 221897
rect 22561 221869 22589 221897
rect 22623 221869 22651 221897
rect 22437 221807 22465 221835
rect 22499 221807 22527 221835
rect 22561 221807 22589 221835
rect 22623 221807 22651 221835
rect 22437 221745 22465 221773
rect 22499 221745 22527 221773
rect 22561 221745 22589 221773
rect 22623 221745 22651 221773
rect 24939 221931 24967 221959
rect 25001 221931 25029 221959
rect 24939 221869 24967 221897
rect 25001 221869 25029 221897
rect 24939 221807 24967 221835
rect 25001 221807 25029 221835
rect 24939 221745 24967 221773
rect 25001 221745 25029 221773
rect 29577 218931 29605 218959
rect 29639 218931 29667 218959
rect 29701 218931 29729 218959
rect 29763 218931 29791 218959
rect 29577 218869 29605 218897
rect 29639 218869 29667 218897
rect 29701 218869 29729 218897
rect 29763 218869 29791 218897
rect 29577 218807 29605 218835
rect 29639 218807 29667 218835
rect 29701 218807 29729 218835
rect 29763 218807 29791 218835
rect 29577 218745 29605 218773
rect 29639 218745 29667 218773
rect 29701 218745 29729 218773
rect 29763 218745 29791 218773
rect 22437 212931 22465 212959
rect 22499 212931 22527 212959
rect 22561 212931 22589 212959
rect 22623 212931 22651 212959
rect 22437 212869 22465 212897
rect 22499 212869 22527 212897
rect 22561 212869 22589 212897
rect 22623 212869 22651 212897
rect 22437 212807 22465 212835
rect 22499 212807 22527 212835
rect 22561 212807 22589 212835
rect 22623 212807 22651 212835
rect 22437 212745 22465 212773
rect 22499 212745 22527 212773
rect 22561 212745 22589 212773
rect 22623 212745 22651 212773
rect 24939 212931 24967 212959
rect 25001 212931 25029 212959
rect 24939 212869 24967 212897
rect 25001 212869 25029 212897
rect 24939 212807 24967 212835
rect 25001 212807 25029 212835
rect 24939 212745 24967 212773
rect 25001 212745 25029 212773
rect 29577 209931 29605 209959
rect 29639 209931 29667 209959
rect 29701 209931 29729 209959
rect 29763 209931 29791 209959
rect 29577 209869 29605 209897
rect 29639 209869 29667 209897
rect 29701 209869 29729 209897
rect 29763 209869 29791 209897
rect 29577 209807 29605 209835
rect 29639 209807 29667 209835
rect 29701 209807 29729 209835
rect 29763 209807 29791 209835
rect 29577 209745 29605 209773
rect 29639 209745 29667 209773
rect 29701 209745 29729 209773
rect 29763 209745 29791 209773
rect 22437 203931 22465 203959
rect 22499 203931 22527 203959
rect 22561 203931 22589 203959
rect 22623 203931 22651 203959
rect 22437 203869 22465 203897
rect 22499 203869 22527 203897
rect 22561 203869 22589 203897
rect 22623 203869 22651 203897
rect 22437 203807 22465 203835
rect 22499 203807 22527 203835
rect 22561 203807 22589 203835
rect 22623 203807 22651 203835
rect 22437 203745 22465 203773
rect 22499 203745 22527 203773
rect 22561 203745 22589 203773
rect 22623 203745 22651 203773
rect 24939 203931 24967 203959
rect 25001 203931 25029 203959
rect 24939 203869 24967 203897
rect 25001 203869 25029 203897
rect 24939 203807 24967 203835
rect 25001 203807 25029 203835
rect 24939 203745 24967 203773
rect 25001 203745 25029 203773
rect 29577 200931 29605 200959
rect 29639 200931 29667 200959
rect 29701 200931 29729 200959
rect 29763 200931 29791 200959
rect 29577 200869 29605 200897
rect 29639 200869 29667 200897
rect 29701 200869 29729 200897
rect 29763 200869 29791 200897
rect 29577 200807 29605 200835
rect 29639 200807 29667 200835
rect 29701 200807 29729 200835
rect 29763 200807 29791 200835
rect 29577 200745 29605 200773
rect 29639 200745 29667 200773
rect 29701 200745 29729 200773
rect 29763 200745 29791 200773
rect 22437 194931 22465 194959
rect 22499 194931 22527 194959
rect 22561 194931 22589 194959
rect 22623 194931 22651 194959
rect 22437 194869 22465 194897
rect 22499 194869 22527 194897
rect 22561 194869 22589 194897
rect 22623 194869 22651 194897
rect 22437 194807 22465 194835
rect 22499 194807 22527 194835
rect 22561 194807 22589 194835
rect 22623 194807 22651 194835
rect 22437 194745 22465 194773
rect 22499 194745 22527 194773
rect 22561 194745 22589 194773
rect 22623 194745 22651 194773
rect 24939 194931 24967 194959
rect 25001 194931 25029 194959
rect 24939 194869 24967 194897
rect 25001 194869 25029 194897
rect 24939 194807 24967 194835
rect 25001 194807 25029 194835
rect 24939 194745 24967 194773
rect 25001 194745 25029 194773
rect 29577 191931 29605 191959
rect 29639 191931 29667 191959
rect 29701 191931 29729 191959
rect 29763 191931 29791 191959
rect 29577 191869 29605 191897
rect 29639 191869 29667 191897
rect 29701 191869 29729 191897
rect 29763 191869 29791 191897
rect 29577 191807 29605 191835
rect 29639 191807 29667 191835
rect 29701 191807 29729 191835
rect 29763 191807 29791 191835
rect 29577 191745 29605 191773
rect 29639 191745 29667 191773
rect 29701 191745 29729 191773
rect 29763 191745 29791 191773
rect 22437 185931 22465 185959
rect 22499 185931 22527 185959
rect 22561 185931 22589 185959
rect 22623 185931 22651 185959
rect 22437 185869 22465 185897
rect 22499 185869 22527 185897
rect 22561 185869 22589 185897
rect 22623 185869 22651 185897
rect 22437 185807 22465 185835
rect 22499 185807 22527 185835
rect 22561 185807 22589 185835
rect 22623 185807 22651 185835
rect 22437 185745 22465 185773
rect 22499 185745 22527 185773
rect 22561 185745 22589 185773
rect 22623 185745 22651 185773
rect 24939 185931 24967 185959
rect 25001 185931 25029 185959
rect 24939 185869 24967 185897
rect 25001 185869 25029 185897
rect 24939 185807 24967 185835
rect 25001 185807 25029 185835
rect 24939 185745 24967 185773
rect 25001 185745 25029 185773
rect 29577 182931 29605 182959
rect 29639 182931 29667 182959
rect 29701 182931 29729 182959
rect 29763 182931 29791 182959
rect 29577 182869 29605 182897
rect 29639 182869 29667 182897
rect 29701 182869 29729 182897
rect 29763 182869 29791 182897
rect 29577 182807 29605 182835
rect 29639 182807 29667 182835
rect 29701 182807 29729 182835
rect 29763 182807 29791 182835
rect 29577 182745 29605 182773
rect 29639 182745 29667 182773
rect 29701 182745 29729 182773
rect 29763 182745 29791 182773
rect 22437 176931 22465 176959
rect 22499 176931 22527 176959
rect 22561 176931 22589 176959
rect 22623 176931 22651 176959
rect 22437 176869 22465 176897
rect 22499 176869 22527 176897
rect 22561 176869 22589 176897
rect 22623 176869 22651 176897
rect 22437 176807 22465 176835
rect 22499 176807 22527 176835
rect 22561 176807 22589 176835
rect 22623 176807 22651 176835
rect 22437 176745 22465 176773
rect 22499 176745 22527 176773
rect 22561 176745 22589 176773
rect 22623 176745 22651 176773
rect 24939 176931 24967 176959
rect 25001 176931 25029 176959
rect 24939 176869 24967 176897
rect 25001 176869 25029 176897
rect 24939 176807 24967 176835
rect 25001 176807 25029 176835
rect 24939 176745 24967 176773
rect 25001 176745 25029 176773
rect 29577 173931 29605 173959
rect 29639 173931 29667 173959
rect 29701 173931 29729 173959
rect 29763 173931 29791 173959
rect 29577 173869 29605 173897
rect 29639 173869 29667 173897
rect 29701 173869 29729 173897
rect 29763 173869 29791 173897
rect 29577 173807 29605 173835
rect 29639 173807 29667 173835
rect 29701 173807 29729 173835
rect 29763 173807 29791 173835
rect 29577 173745 29605 173773
rect 29639 173745 29667 173773
rect 29701 173745 29729 173773
rect 29763 173745 29791 173773
rect 22437 167931 22465 167959
rect 22499 167931 22527 167959
rect 22561 167931 22589 167959
rect 22623 167931 22651 167959
rect 22437 167869 22465 167897
rect 22499 167869 22527 167897
rect 22561 167869 22589 167897
rect 22623 167869 22651 167897
rect 22437 167807 22465 167835
rect 22499 167807 22527 167835
rect 22561 167807 22589 167835
rect 22623 167807 22651 167835
rect 22437 167745 22465 167773
rect 22499 167745 22527 167773
rect 22561 167745 22589 167773
rect 22623 167745 22651 167773
rect 24939 167931 24967 167959
rect 25001 167931 25029 167959
rect 24939 167869 24967 167897
rect 25001 167869 25029 167897
rect 24939 167807 24967 167835
rect 25001 167807 25029 167835
rect 24939 167745 24967 167773
rect 25001 167745 25029 167773
rect 29577 164931 29605 164959
rect 29639 164931 29667 164959
rect 29701 164931 29729 164959
rect 29763 164931 29791 164959
rect 29577 164869 29605 164897
rect 29639 164869 29667 164897
rect 29701 164869 29729 164897
rect 29763 164869 29791 164897
rect 29577 164807 29605 164835
rect 29639 164807 29667 164835
rect 29701 164807 29729 164835
rect 29763 164807 29791 164835
rect 29577 164745 29605 164773
rect 29639 164745 29667 164773
rect 29701 164745 29729 164773
rect 29763 164745 29791 164773
rect 22437 158931 22465 158959
rect 22499 158931 22527 158959
rect 22561 158931 22589 158959
rect 22623 158931 22651 158959
rect 22437 158869 22465 158897
rect 22499 158869 22527 158897
rect 22561 158869 22589 158897
rect 22623 158869 22651 158897
rect 22437 158807 22465 158835
rect 22499 158807 22527 158835
rect 22561 158807 22589 158835
rect 22623 158807 22651 158835
rect 22437 158745 22465 158773
rect 22499 158745 22527 158773
rect 22561 158745 22589 158773
rect 22623 158745 22651 158773
rect 24939 158931 24967 158959
rect 25001 158931 25029 158959
rect 24939 158869 24967 158897
rect 25001 158869 25029 158897
rect 24939 158807 24967 158835
rect 25001 158807 25029 158835
rect 24939 158745 24967 158773
rect 25001 158745 25029 158773
rect 29577 155931 29605 155959
rect 29639 155931 29667 155959
rect 29701 155931 29729 155959
rect 29763 155931 29791 155959
rect 29577 155869 29605 155897
rect 29639 155869 29667 155897
rect 29701 155869 29729 155897
rect 29763 155869 29791 155897
rect 29577 155807 29605 155835
rect 29639 155807 29667 155835
rect 29701 155807 29729 155835
rect 29763 155807 29791 155835
rect 29577 155745 29605 155773
rect 29639 155745 29667 155773
rect 29701 155745 29729 155773
rect 29763 155745 29791 155773
rect 22437 149931 22465 149959
rect 22499 149931 22527 149959
rect 22561 149931 22589 149959
rect 22623 149931 22651 149959
rect 22437 149869 22465 149897
rect 22499 149869 22527 149897
rect 22561 149869 22589 149897
rect 22623 149869 22651 149897
rect 22437 149807 22465 149835
rect 22499 149807 22527 149835
rect 22561 149807 22589 149835
rect 22623 149807 22651 149835
rect 22437 149745 22465 149773
rect 22499 149745 22527 149773
rect 22561 149745 22589 149773
rect 22623 149745 22651 149773
rect 24939 149931 24967 149959
rect 25001 149931 25029 149959
rect 24939 149869 24967 149897
rect 25001 149869 25029 149897
rect 24939 149807 24967 149835
rect 25001 149807 25029 149835
rect 24939 149745 24967 149773
rect 25001 149745 25029 149773
rect 29577 146931 29605 146959
rect 29639 146931 29667 146959
rect 29701 146931 29729 146959
rect 29763 146931 29791 146959
rect 29577 146869 29605 146897
rect 29639 146869 29667 146897
rect 29701 146869 29729 146897
rect 29763 146869 29791 146897
rect 29577 146807 29605 146835
rect 29639 146807 29667 146835
rect 29701 146807 29729 146835
rect 29763 146807 29791 146835
rect 29577 146745 29605 146773
rect 29639 146745 29667 146773
rect 29701 146745 29729 146773
rect 29763 146745 29791 146773
rect 22437 140931 22465 140959
rect 22499 140931 22527 140959
rect 22561 140931 22589 140959
rect 22623 140931 22651 140959
rect 22437 140869 22465 140897
rect 22499 140869 22527 140897
rect 22561 140869 22589 140897
rect 22623 140869 22651 140897
rect 22437 140807 22465 140835
rect 22499 140807 22527 140835
rect 22561 140807 22589 140835
rect 22623 140807 22651 140835
rect 22437 140745 22465 140773
rect 22499 140745 22527 140773
rect 22561 140745 22589 140773
rect 22623 140745 22651 140773
rect 24939 140931 24967 140959
rect 25001 140931 25029 140959
rect 24939 140869 24967 140897
rect 25001 140869 25029 140897
rect 24939 140807 24967 140835
rect 25001 140807 25029 140835
rect 24939 140745 24967 140773
rect 25001 140745 25029 140773
rect 29577 137931 29605 137959
rect 29639 137931 29667 137959
rect 29701 137931 29729 137959
rect 29763 137931 29791 137959
rect 29577 137869 29605 137897
rect 29639 137869 29667 137897
rect 29701 137869 29729 137897
rect 29763 137869 29791 137897
rect 29577 137807 29605 137835
rect 29639 137807 29667 137835
rect 29701 137807 29729 137835
rect 29763 137807 29791 137835
rect 29577 137745 29605 137773
rect 29639 137745 29667 137773
rect 29701 137745 29729 137773
rect 29763 137745 29791 137773
rect 22437 131931 22465 131959
rect 22499 131931 22527 131959
rect 22561 131931 22589 131959
rect 22623 131931 22651 131959
rect 22437 131869 22465 131897
rect 22499 131869 22527 131897
rect 22561 131869 22589 131897
rect 22623 131869 22651 131897
rect 22437 131807 22465 131835
rect 22499 131807 22527 131835
rect 22561 131807 22589 131835
rect 22623 131807 22651 131835
rect 22437 131745 22465 131773
rect 22499 131745 22527 131773
rect 22561 131745 22589 131773
rect 22623 131745 22651 131773
rect 24939 131931 24967 131959
rect 25001 131931 25029 131959
rect 24939 131869 24967 131897
rect 25001 131869 25029 131897
rect 24939 131807 24967 131835
rect 25001 131807 25029 131835
rect 24939 131745 24967 131773
rect 25001 131745 25029 131773
rect 29577 128931 29605 128959
rect 29639 128931 29667 128959
rect 29701 128931 29729 128959
rect 29763 128931 29791 128959
rect 29577 128869 29605 128897
rect 29639 128869 29667 128897
rect 29701 128869 29729 128897
rect 29763 128869 29791 128897
rect 29577 128807 29605 128835
rect 29639 128807 29667 128835
rect 29701 128807 29729 128835
rect 29763 128807 29791 128835
rect 29577 128745 29605 128773
rect 29639 128745 29667 128773
rect 29701 128745 29729 128773
rect 29763 128745 29791 128773
rect 22437 122931 22465 122959
rect 22499 122931 22527 122959
rect 22561 122931 22589 122959
rect 22623 122931 22651 122959
rect 22437 122869 22465 122897
rect 22499 122869 22527 122897
rect 22561 122869 22589 122897
rect 22623 122869 22651 122897
rect 22437 122807 22465 122835
rect 22499 122807 22527 122835
rect 22561 122807 22589 122835
rect 22623 122807 22651 122835
rect 22437 122745 22465 122773
rect 22499 122745 22527 122773
rect 22561 122745 22589 122773
rect 22623 122745 22651 122773
rect 24939 122931 24967 122959
rect 25001 122931 25029 122959
rect 24939 122869 24967 122897
rect 25001 122869 25029 122897
rect 24939 122807 24967 122835
rect 25001 122807 25029 122835
rect 24939 122745 24967 122773
rect 25001 122745 25029 122773
rect 29577 119931 29605 119959
rect 29639 119931 29667 119959
rect 29701 119931 29729 119959
rect 29763 119931 29791 119959
rect 29577 119869 29605 119897
rect 29639 119869 29667 119897
rect 29701 119869 29729 119897
rect 29763 119869 29791 119897
rect 29577 119807 29605 119835
rect 29639 119807 29667 119835
rect 29701 119807 29729 119835
rect 29763 119807 29791 119835
rect 29577 119745 29605 119773
rect 29639 119745 29667 119773
rect 29701 119745 29729 119773
rect 29763 119745 29791 119773
rect 22437 113931 22465 113959
rect 22499 113931 22527 113959
rect 22561 113931 22589 113959
rect 22623 113931 22651 113959
rect 22437 113869 22465 113897
rect 22499 113869 22527 113897
rect 22561 113869 22589 113897
rect 22623 113869 22651 113897
rect 22437 113807 22465 113835
rect 22499 113807 22527 113835
rect 22561 113807 22589 113835
rect 22623 113807 22651 113835
rect 22437 113745 22465 113773
rect 22499 113745 22527 113773
rect 22561 113745 22589 113773
rect 22623 113745 22651 113773
rect 24939 113931 24967 113959
rect 25001 113931 25029 113959
rect 24939 113869 24967 113897
rect 25001 113869 25029 113897
rect 24939 113807 24967 113835
rect 25001 113807 25029 113835
rect 24939 113745 24967 113773
rect 25001 113745 25029 113773
rect 29577 110931 29605 110959
rect 29639 110931 29667 110959
rect 29701 110931 29729 110959
rect 29763 110931 29791 110959
rect 29577 110869 29605 110897
rect 29639 110869 29667 110897
rect 29701 110869 29729 110897
rect 29763 110869 29791 110897
rect 29577 110807 29605 110835
rect 29639 110807 29667 110835
rect 29701 110807 29729 110835
rect 29763 110807 29791 110835
rect 29577 110745 29605 110773
rect 29639 110745 29667 110773
rect 29701 110745 29729 110773
rect 29763 110745 29791 110773
rect 22437 104931 22465 104959
rect 22499 104931 22527 104959
rect 22561 104931 22589 104959
rect 22623 104931 22651 104959
rect 22437 104869 22465 104897
rect 22499 104869 22527 104897
rect 22561 104869 22589 104897
rect 22623 104869 22651 104897
rect 22437 104807 22465 104835
rect 22499 104807 22527 104835
rect 22561 104807 22589 104835
rect 22623 104807 22651 104835
rect 22437 104745 22465 104773
rect 22499 104745 22527 104773
rect 22561 104745 22589 104773
rect 22623 104745 22651 104773
rect 24939 104931 24967 104959
rect 25001 104931 25029 104959
rect 24939 104869 24967 104897
rect 25001 104869 25029 104897
rect 24939 104807 24967 104835
rect 25001 104807 25029 104835
rect 24939 104745 24967 104773
rect 25001 104745 25029 104773
rect 29577 101931 29605 101959
rect 29639 101931 29667 101959
rect 29701 101931 29729 101959
rect 29763 101931 29791 101959
rect 29577 101869 29605 101897
rect 29639 101869 29667 101897
rect 29701 101869 29729 101897
rect 29763 101869 29791 101897
rect 29577 101807 29605 101835
rect 29639 101807 29667 101835
rect 29701 101807 29729 101835
rect 29763 101807 29791 101835
rect 29577 101745 29605 101773
rect 29639 101745 29667 101773
rect 29701 101745 29729 101773
rect 29763 101745 29791 101773
rect 22437 95931 22465 95959
rect 22499 95931 22527 95959
rect 22561 95931 22589 95959
rect 22623 95931 22651 95959
rect 22437 95869 22465 95897
rect 22499 95869 22527 95897
rect 22561 95869 22589 95897
rect 22623 95869 22651 95897
rect 22437 95807 22465 95835
rect 22499 95807 22527 95835
rect 22561 95807 22589 95835
rect 22623 95807 22651 95835
rect 22437 95745 22465 95773
rect 22499 95745 22527 95773
rect 22561 95745 22589 95773
rect 22623 95745 22651 95773
rect 24939 95931 24967 95959
rect 25001 95931 25029 95959
rect 24939 95869 24967 95897
rect 25001 95869 25029 95897
rect 24939 95807 24967 95835
rect 25001 95807 25029 95835
rect 24939 95745 24967 95773
rect 25001 95745 25029 95773
rect 29577 92931 29605 92959
rect 29639 92931 29667 92959
rect 29701 92931 29729 92959
rect 29763 92931 29791 92959
rect 29577 92869 29605 92897
rect 29639 92869 29667 92897
rect 29701 92869 29729 92897
rect 29763 92869 29791 92897
rect 29577 92807 29605 92835
rect 29639 92807 29667 92835
rect 29701 92807 29729 92835
rect 29763 92807 29791 92835
rect 29577 92745 29605 92773
rect 29639 92745 29667 92773
rect 29701 92745 29729 92773
rect 29763 92745 29791 92773
rect 22437 86931 22465 86959
rect 22499 86931 22527 86959
rect 22561 86931 22589 86959
rect 22623 86931 22651 86959
rect 22437 86869 22465 86897
rect 22499 86869 22527 86897
rect 22561 86869 22589 86897
rect 22623 86869 22651 86897
rect 22437 86807 22465 86835
rect 22499 86807 22527 86835
rect 22561 86807 22589 86835
rect 22623 86807 22651 86835
rect 22437 86745 22465 86773
rect 22499 86745 22527 86773
rect 22561 86745 22589 86773
rect 22623 86745 22651 86773
rect 24939 86931 24967 86959
rect 25001 86931 25029 86959
rect 24939 86869 24967 86897
rect 25001 86869 25029 86897
rect 24939 86807 24967 86835
rect 25001 86807 25029 86835
rect 24939 86745 24967 86773
rect 25001 86745 25029 86773
rect 29577 83931 29605 83959
rect 29639 83931 29667 83959
rect 29701 83931 29729 83959
rect 29763 83931 29791 83959
rect 29577 83869 29605 83897
rect 29639 83869 29667 83897
rect 29701 83869 29729 83897
rect 29763 83869 29791 83897
rect 29577 83807 29605 83835
rect 29639 83807 29667 83835
rect 29701 83807 29729 83835
rect 29763 83807 29791 83835
rect 29577 83745 29605 83773
rect 29639 83745 29667 83773
rect 29701 83745 29729 83773
rect 29763 83745 29791 83773
rect 22437 77931 22465 77959
rect 22499 77931 22527 77959
rect 22561 77931 22589 77959
rect 22623 77931 22651 77959
rect 22437 77869 22465 77897
rect 22499 77869 22527 77897
rect 22561 77869 22589 77897
rect 22623 77869 22651 77897
rect 22437 77807 22465 77835
rect 22499 77807 22527 77835
rect 22561 77807 22589 77835
rect 22623 77807 22651 77835
rect 22437 77745 22465 77773
rect 22499 77745 22527 77773
rect 22561 77745 22589 77773
rect 22623 77745 22651 77773
rect 24939 77931 24967 77959
rect 25001 77931 25029 77959
rect 24939 77869 24967 77897
rect 25001 77869 25029 77897
rect 24939 77807 24967 77835
rect 25001 77807 25029 77835
rect 24939 77745 24967 77773
rect 25001 77745 25029 77773
rect 29577 74931 29605 74959
rect 29639 74931 29667 74959
rect 29701 74931 29729 74959
rect 29763 74931 29791 74959
rect 29577 74869 29605 74897
rect 29639 74869 29667 74897
rect 29701 74869 29729 74897
rect 29763 74869 29791 74897
rect 29577 74807 29605 74835
rect 29639 74807 29667 74835
rect 29701 74807 29729 74835
rect 29763 74807 29791 74835
rect 29577 74745 29605 74773
rect 29639 74745 29667 74773
rect 29701 74745 29729 74773
rect 29763 74745 29791 74773
rect 22437 68931 22465 68959
rect 22499 68931 22527 68959
rect 22561 68931 22589 68959
rect 22623 68931 22651 68959
rect 22437 68869 22465 68897
rect 22499 68869 22527 68897
rect 22561 68869 22589 68897
rect 22623 68869 22651 68897
rect 22437 68807 22465 68835
rect 22499 68807 22527 68835
rect 22561 68807 22589 68835
rect 22623 68807 22651 68835
rect 22437 68745 22465 68773
rect 22499 68745 22527 68773
rect 22561 68745 22589 68773
rect 22623 68745 22651 68773
rect 24939 68931 24967 68959
rect 25001 68931 25029 68959
rect 24939 68869 24967 68897
rect 25001 68869 25029 68897
rect 24939 68807 24967 68835
rect 25001 68807 25029 68835
rect 24939 68745 24967 68773
rect 25001 68745 25029 68773
rect 29577 65931 29605 65959
rect 29639 65931 29667 65959
rect 29701 65931 29729 65959
rect 29763 65931 29791 65959
rect 29577 65869 29605 65897
rect 29639 65869 29667 65897
rect 29701 65869 29729 65897
rect 29763 65869 29791 65897
rect 29577 65807 29605 65835
rect 29639 65807 29667 65835
rect 29701 65807 29729 65835
rect 29763 65807 29791 65835
rect 29577 65745 29605 65773
rect 29639 65745 29667 65773
rect 29701 65745 29729 65773
rect 29763 65745 29791 65773
rect 22437 59931 22465 59959
rect 22499 59931 22527 59959
rect 22561 59931 22589 59959
rect 22623 59931 22651 59959
rect 22437 59869 22465 59897
rect 22499 59869 22527 59897
rect 22561 59869 22589 59897
rect 22623 59869 22651 59897
rect 22437 59807 22465 59835
rect 22499 59807 22527 59835
rect 22561 59807 22589 59835
rect 22623 59807 22651 59835
rect 22437 59745 22465 59773
rect 22499 59745 22527 59773
rect 22561 59745 22589 59773
rect 22623 59745 22651 59773
rect 24939 59931 24967 59959
rect 25001 59931 25029 59959
rect 24939 59869 24967 59897
rect 25001 59869 25029 59897
rect 24939 59807 24967 59835
rect 25001 59807 25029 59835
rect 24939 59745 24967 59773
rect 25001 59745 25029 59773
rect 29577 56931 29605 56959
rect 29639 56931 29667 56959
rect 29701 56931 29729 56959
rect 29763 56931 29791 56959
rect 29577 56869 29605 56897
rect 29639 56869 29667 56897
rect 29701 56869 29729 56897
rect 29763 56869 29791 56897
rect 29577 56807 29605 56835
rect 29639 56807 29667 56835
rect 29701 56807 29729 56835
rect 29763 56807 29791 56835
rect 29577 56745 29605 56773
rect 29639 56745 29667 56773
rect 29701 56745 29729 56773
rect 29763 56745 29791 56773
rect 22437 50931 22465 50959
rect 22499 50931 22527 50959
rect 22561 50931 22589 50959
rect 22623 50931 22651 50959
rect 22437 50869 22465 50897
rect 22499 50869 22527 50897
rect 22561 50869 22589 50897
rect 22623 50869 22651 50897
rect 22437 50807 22465 50835
rect 22499 50807 22527 50835
rect 22561 50807 22589 50835
rect 22623 50807 22651 50835
rect 22437 50745 22465 50773
rect 22499 50745 22527 50773
rect 22561 50745 22589 50773
rect 22623 50745 22651 50773
rect 24939 50931 24967 50959
rect 25001 50931 25029 50959
rect 24939 50869 24967 50897
rect 25001 50869 25029 50897
rect 24939 50807 24967 50835
rect 25001 50807 25029 50835
rect 24939 50745 24967 50773
rect 25001 50745 25029 50773
rect 29577 47931 29605 47959
rect 29639 47931 29667 47959
rect 29701 47931 29729 47959
rect 29763 47931 29791 47959
rect 29577 47869 29605 47897
rect 29639 47869 29667 47897
rect 29701 47869 29729 47897
rect 29763 47869 29791 47897
rect 29577 47807 29605 47835
rect 29639 47807 29667 47835
rect 29701 47807 29729 47835
rect 29763 47807 29791 47835
rect 29577 47745 29605 47773
rect 29639 47745 29667 47773
rect 29701 47745 29729 47773
rect 29763 47745 29791 47773
rect 22437 41931 22465 41959
rect 22499 41931 22527 41959
rect 22561 41931 22589 41959
rect 22623 41931 22651 41959
rect 22437 41869 22465 41897
rect 22499 41869 22527 41897
rect 22561 41869 22589 41897
rect 22623 41869 22651 41897
rect 22437 41807 22465 41835
rect 22499 41807 22527 41835
rect 22561 41807 22589 41835
rect 22623 41807 22651 41835
rect 22437 41745 22465 41773
rect 22499 41745 22527 41773
rect 22561 41745 22589 41773
rect 22623 41745 22651 41773
rect 24939 41931 24967 41959
rect 25001 41931 25029 41959
rect 24939 41869 24967 41897
rect 25001 41869 25029 41897
rect 24939 41807 24967 41835
rect 25001 41807 25029 41835
rect 24939 41745 24967 41773
rect 25001 41745 25029 41773
rect 29577 38931 29605 38959
rect 29639 38931 29667 38959
rect 29701 38931 29729 38959
rect 29763 38931 29791 38959
rect 29577 38869 29605 38897
rect 29639 38869 29667 38897
rect 29701 38869 29729 38897
rect 29763 38869 29791 38897
rect 29577 38807 29605 38835
rect 29639 38807 29667 38835
rect 29701 38807 29729 38835
rect 29763 38807 29791 38835
rect 29577 38745 29605 38773
rect 29639 38745 29667 38773
rect 29701 38745 29729 38773
rect 29763 38745 29791 38773
rect 22437 32931 22465 32959
rect 22499 32931 22527 32959
rect 22561 32931 22589 32959
rect 22623 32931 22651 32959
rect 22437 32869 22465 32897
rect 22499 32869 22527 32897
rect 22561 32869 22589 32897
rect 22623 32869 22651 32897
rect 22437 32807 22465 32835
rect 22499 32807 22527 32835
rect 22561 32807 22589 32835
rect 22623 32807 22651 32835
rect 22437 32745 22465 32773
rect 22499 32745 22527 32773
rect 22561 32745 22589 32773
rect 22623 32745 22651 32773
rect 24939 32931 24967 32959
rect 25001 32931 25029 32959
rect 24939 32869 24967 32897
rect 25001 32869 25029 32897
rect 24939 32807 24967 32835
rect 25001 32807 25029 32835
rect 24939 32745 24967 32773
rect 25001 32745 25029 32773
rect 29577 29931 29605 29959
rect 29639 29931 29667 29959
rect 29701 29931 29729 29959
rect 29763 29931 29791 29959
rect 29577 29869 29605 29897
rect 29639 29869 29667 29897
rect 29701 29869 29729 29897
rect 29763 29869 29791 29897
rect 29577 29807 29605 29835
rect 29639 29807 29667 29835
rect 29701 29807 29729 29835
rect 29763 29807 29791 29835
rect 29577 29745 29605 29773
rect 29639 29745 29667 29773
rect 29701 29745 29729 29773
rect 29763 29745 29791 29773
rect 22437 23931 22465 23959
rect 22499 23931 22527 23959
rect 22561 23931 22589 23959
rect 22623 23931 22651 23959
rect 22437 23869 22465 23897
rect 22499 23869 22527 23897
rect 22561 23869 22589 23897
rect 22623 23869 22651 23897
rect 22437 23807 22465 23835
rect 22499 23807 22527 23835
rect 22561 23807 22589 23835
rect 22623 23807 22651 23835
rect 22437 23745 22465 23773
rect 22499 23745 22527 23773
rect 22561 23745 22589 23773
rect 22623 23745 22651 23773
rect 24939 23931 24967 23959
rect 25001 23931 25029 23959
rect 24939 23869 24967 23897
rect 25001 23869 25029 23897
rect 24939 23807 24967 23835
rect 25001 23807 25029 23835
rect 24939 23745 24967 23773
rect 25001 23745 25029 23773
rect 22437 14931 22465 14959
rect 22499 14931 22527 14959
rect 22561 14931 22589 14959
rect 22623 14931 22651 14959
rect 22437 14869 22465 14897
rect 22499 14869 22527 14897
rect 22561 14869 22589 14897
rect 22623 14869 22651 14897
rect 22437 14807 22465 14835
rect 22499 14807 22527 14835
rect 22561 14807 22589 14835
rect 22623 14807 22651 14835
rect 22437 14745 22465 14773
rect 22499 14745 22527 14773
rect 22561 14745 22589 14773
rect 22623 14745 22651 14773
rect 22437 5931 22465 5959
rect 22499 5931 22527 5959
rect 22561 5931 22589 5959
rect 22623 5931 22651 5959
rect 22437 5869 22465 5897
rect 22499 5869 22527 5897
rect 22561 5869 22589 5897
rect 22623 5869 22651 5897
rect 22437 5807 22465 5835
rect 22499 5807 22527 5835
rect 22561 5807 22589 5835
rect 22623 5807 22651 5835
rect 22437 5745 22465 5773
rect 22499 5745 22527 5773
rect 22561 5745 22589 5773
rect 22623 5745 22651 5773
rect 22437 396 22465 424
rect 22499 396 22527 424
rect 22561 396 22589 424
rect 22623 396 22651 424
rect 22437 334 22465 362
rect 22499 334 22527 362
rect 22561 334 22589 362
rect 22623 334 22651 362
rect 22437 272 22465 300
rect 22499 272 22527 300
rect 22561 272 22589 300
rect 22623 272 22651 300
rect 22437 210 22465 238
rect 22499 210 22527 238
rect 22561 210 22589 238
rect 22623 210 22651 238
rect 29577 20931 29605 20959
rect 29639 20931 29667 20959
rect 29701 20931 29729 20959
rect 29763 20931 29791 20959
rect 29577 20869 29605 20897
rect 29639 20869 29667 20897
rect 29701 20869 29729 20897
rect 29763 20869 29791 20897
rect 29577 20807 29605 20835
rect 29639 20807 29667 20835
rect 29701 20807 29729 20835
rect 29763 20807 29791 20835
rect 29577 20745 29605 20773
rect 29639 20745 29667 20773
rect 29701 20745 29729 20773
rect 29763 20745 29791 20773
rect 29577 11931 29605 11959
rect 29639 11931 29667 11959
rect 29701 11931 29729 11959
rect 29763 11931 29791 11959
rect 29577 11869 29605 11897
rect 29639 11869 29667 11897
rect 29701 11869 29729 11897
rect 29763 11869 29791 11897
rect 29577 11807 29605 11835
rect 29639 11807 29667 11835
rect 29701 11807 29729 11835
rect 29763 11807 29791 11835
rect 29577 11745 29605 11773
rect 29639 11745 29667 11773
rect 29701 11745 29729 11773
rect 29763 11745 29791 11773
rect 29577 2931 29605 2959
rect 29639 2931 29667 2959
rect 29701 2931 29729 2959
rect 29763 2931 29791 2959
rect 29577 2869 29605 2897
rect 29639 2869 29667 2897
rect 29701 2869 29729 2897
rect 29763 2869 29791 2897
rect 29577 2807 29605 2835
rect 29639 2807 29667 2835
rect 29701 2807 29729 2835
rect 29763 2807 29791 2835
rect 29577 2745 29605 2773
rect 29639 2745 29667 2773
rect 29701 2745 29729 2773
rect 29763 2745 29791 2773
rect 29577 876 29605 904
rect 29639 876 29667 904
rect 29701 876 29729 904
rect 29763 876 29791 904
rect 29577 814 29605 842
rect 29639 814 29667 842
rect 29701 814 29729 842
rect 29763 814 29791 842
rect 29577 752 29605 780
rect 29639 752 29667 780
rect 29701 752 29729 780
rect 29763 752 29791 780
rect 29577 690 29605 718
rect 29639 690 29667 718
rect 29701 690 29729 718
rect 29763 690 29791 718
rect 31437 299642 31465 299670
rect 31499 299642 31527 299670
rect 31561 299642 31589 299670
rect 31623 299642 31651 299670
rect 31437 299580 31465 299608
rect 31499 299580 31527 299608
rect 31561 299580 31589 299608
rect 31623 299580 31651 299608
rect 31437 299518 31465 299546
rect 31499 299518 31527 299546
rect 31561 299518 31589 299546
rect 31623 299518 31651 299546
rect 31437 299456 31465 299484
rect 31499 299456 31527 299484
rect 31561 299456 31589 299484
rect 31623 299456 31651 299484
rect 31437 293931 31465 293959
rect 31499 293931 31527 293959
rect 31561 293931 31589 293959
rect 31623 293931 31651 293959
rect 31437 293869 31465 293897
rect 31499 293869 31527 293897
rect 31561 293869 31589 293897
rect 31623 293869 31651 293897
rect 31437 293807 31465 293835
rect 31499 293807 31527 293835
rect 31561 293807 31589 293835
rect 31623 293807 31651 293835
rect 31437 293745 31465 293773
rect 31499 293745 31527 293773
rect 31561 293745 31589 293773
rect 31623 293745 31651 293773
rect 31437 284931 31465 284959
rect 31499 284931 31527 284959
rect 31561 284931 31589 284959
rect 31623 284931 31651 284959
rect 31437 284869 31465 284897
rect 31499 284869 31527 284897
rect 31561 284869 31589 284897
rect 31623 284869 31651 284897
rect 31437 284807 31465 284835
rect 31499 284807 31527 284835
rect 31561 284807 31589 284835
rect 31623 284807 31651 284835
rect 31437 284745 31465 284773
rect 31499 284745 31527 284773
rect 31561 284745 31589 284773
rect 31623 284745 31651 284773
rect 31437 275931 31465 275959
rect 31499 275931 31527 275959
rect 31561 275931 31589 275959
rect 31623 275931 31651 275959
rect 31437 275869 31465 275897
rect 31499 275869 31527 275897
rect 31561 275869 31589 275897
rect 31623 275869 31651 275897
rect 31437 275807 31465 275835
rect 31499 275807 31527 275835
rect 31561 275807 31589 275835
rect 31623 275807 31651 275835
rect 31437 275745 31465 275773
rect 31499 275745 31527 275773
rect 31561 275745 31589 275773
rect 31623 275745 31651 275773
rect 31437 266931 31465 266959
rect 31499 266931 31527 266959
rect 31561 266931 31589 266959
rect 31623 266931 31651 266959
rect 31437 266869 31465 266897
rect 31499 266869 31527 266897
rect 31561 266869 31589 266897
rect 31623 266869 31651 266897
rect 31437 266807 31465 266835
rect 31499 266807 31527 266835
rect 31561 266807 31589 266835
rect 31623 266807 31651 266835
rect 31437 266745 31465 266773
rect 31499 266745 31527 266773
rect 31561 266745 31589 266773
rect 31623 266745 31651 266773
rect 31437 257931 31465 257959
rect 31499 257931 31527 257959
rect 31561 257931 31589 257959
rect 31623 257931 31651 257959
rect 31437 257869 31465 257897
rect 31499 257869 31527 257897
rect 31561 257869 31589 257897
rect 31623 257869 31651 257897
rect 31437 257807 31465 257835
rect 31499 257807 31527 257835
rect 31561 257807 31589 257835
rect 31623 257807 31651 257835
rect 31437 257745 31465 257773
rect 31499 257745 31527 257773
rect 31561 257745 31589 257773
rect 31623 257745 31651 257773
rect 38577 299162 38605 299190
rect 38639 299162 38667 299190
rect 38701 299162 38729 299190
rect 38763 299162 38791 299190
rect 38577 299100 38605 299128
rect 38639 299100 38667 299128
rect 38701 299100 38729 299128
rect 38763 299100 38791 299128
rect 38577 299038 38605 299066
rect 38639 299038 38667 299066
rect 38701 299038 38729 299066
rect 38763 299038 38791 299066
rect 38577 298976 38605 299004
rect 38639 298976 38667 299004
rect 38701 298976 38729 299004
rect 38763 298976 38791 299004
rect 38577 290931 38605 290959
rect 38639 290931 38667 290959
rect 38701 290931 38729 290959
rect 38763 290931 38791 290959
rect 38577 290869 38605 290897
rect 38639 290869 38667 290897
rect 38701 290869 38729 290897
rect 38763 290869 38791 290897
rect 38577 290807 38605 290835
rect 38639 290807 38667 290835
rect 38701 290807 38729 290835
rect 38763 290807 38791 290835
rect 38577 290745 38605 290773
rect 38639 290745 38667 290773
rect 38701 290745 38729 290773
rect 38763 290745 38791 290773
rect 38577 281931 38605 281959
rect 38639 281931 38667 281959
rect 38701 281931 38729 281959
rect 38763 281931 38791 281959
rect 38577 281869 38605 281897
rect 38639 281869 38667 281897
rect 38701 281869 38729 281897
rect 38763 281869 38791 281897
rect 38577 281807 38605 281835
rect 38639 281807 38667 281835
rect 38701 281807 38729 281835
rect 38763 281807 38791 281835
rect 38577 281745 38605 281773
rect 38639 281745 38667 281773
rect 38701 281745 38729 281773
rect 38763 281745 38791 281773
rect 38577 272931 38605 272959
rect 38639 272931 38667 272959
rect 38701 272931 38729 272959
rect 38763 272931 38791 272959
rect 38577 272869 38605 272897
rect 38639 272869 38667 272897
rect 38701 272869 38729 272897
rect 38763 272869 38791 272897
rect 38577 272807 38605 272835
rect 38639 272807 38667 272835
rect 38701 272807 38729 272835
rect 38763 272807 38791 272835
rect 38577 272745 38605 272773
rect 38639 272745 38667 272773
rect 38701 272745 38729 272773
rect 38763 272745 38791 272773
rect 38577 263931 38605 263959
rect 38639 263931 38667 263959
rect 38701 263931 38729 263959
rect 38763 263931 38791 263959
rect 38577 263869 38605 263897
rect 38639 263869 38667 263897
rect 38701 263869 38729 263897
rect 38763 263869 38791 263897
rect 38577 263807 38605 263835
rect 38639 263807 38667 263835
rect 38701 263807 38729 263835
rect 38763 263807 38791 263835
rect 38577 263745 38605 263773
rect 38639 263745 38667 263773
rect 38701 263745 38729 263773
rect 38763 263745 38791 263773
rect 38577 254931 38605 254959
rect 38639 254931 38667 254959
rect 38701 254931 38729 254959
rect 38763 254931 38791 254959
rect 38577 254869 38605 254897
rect 38639 254869 38667 254897
rect 38701 254869 38729 254897
rect 38763 254869 38791 254897
rect 38577 254807 38605 254835
rect 38639 254807 38667 254835
rect 38701 254807 38729 254835
rect 38763 254807 38791 254835
rect 38577 254745 38605 254773
rect 38639 254745 38667 254773
rect 38701 254745 38729 254773
rect 38763 254745 38791 254773
rect 40437 299642 40465 299670
rect 40499 299642 40527 299670
rect 40561 299642 40589 299670
rect 40623 299642 40651 299670
rect 40437 299580 40465 299608
rect 40499 299580 40527 299608
rect 40561 299580 40589 299608
rect 40623 299580 40651 299608
rect 40437 299518 40465 299546
rect 40499 299518 40527 299546
rect 40561 299518 40589 299546
rect 40623 299518 40651 299546
rect 40437 299456 40465 299484
rect 40499 299456 40527 299484
rect 40561 299456 40589 299484
rect 40623 299456 40651 299484
rect 40437 293931 40465 293959
rect 40499 293931 40527 293959
rect 40561 293931 40589 293959
rect 40623 293931 40651 293959
rect 40437 293869 40465 293897
rect 40499 293869 40527 293897
rect 40561 293869 40589 293897
rect 40623 293869 40651 293897
rect 40437 293807 40465 293835
rect 40499 293807 40527 293835
rect 40561 293807 40589 293835
rect 40623 293807 40651 293835
rect 40437 293745 40465 293773
rect 40499 293745 40527 293773
rect 40561 293745 40589 293773
rect 40623 293745 40651 293773
rect 40437 284931 40465 284959
rect 40499 284931 40527 284959
rect 40561 284931 40589 284959
rect 40623 284931 40651 284959
rect 40437 284869 40465 284897
rect 40499 284869 40527 284897
rect 40561 284869 40589 284897
rect 40623 284869 40651 284897
rect 40437 284807 40465 284835
rect 40499 284807 40527 284835
rect 40561 284807 40589 284835
rect 40623 284807 40651 284835
rect 40437 284745 40465 284773
rect 40499 284745 40527 284773
rect 40561 284745 40589 284773
rect 40623 284745 40651 284773
rect 40437 275931 40465 275959
rect 40499 275931 40527 275959
rect 40561 275931 40589 275959
rect 40623 275931 40651 275959
rect 40437 275869 40465 275897
rect 40499 275869 40527 275897
rect 40561 275869 40589 275897
rect 40623 275869 40651 275897
rect 40437 275807 40465 275835
rect 40499 275807 40527 275835
rect 40561 275807 40589 275835
rect 40623 275807 40651 275835
rect 40437 275745 40465 275773
rect 40499 275745 40527 275773
rect 40561 275745 40589 275773
rect 40623 275745 40651 275773
rect 40437 266931 40465 266959
rect 40499 266931 40527 266959
rect 40561 266931 40589 266959
rect 40623 266931 40651 266959
rect 40437 266869 40465 266897
rect 40499 266869 40527 266897
rect 40561 266869 40589 266897
rect 40623 266869 40651 266897
rect 40437 266807 40465 266835
rect 40499 266807 40527 266835
rect 40561 266807 40589 266835
rect 40623 266807 40651 266835
rect 40437 266745 40465 266773
rect 40499 266745 40527 266773
rect 40561 266745 40589 266773
rect 40623 266745 40651 266773
rect 40437 257931 40465 257959
rect 40499 257931 40527 257959
rect 40561 257931 40589 257959
rect 40623 257931 40651 257959
rect 40437 257869 40465 257897
rect 40499 257869 40527 257897
rect 40561 257869 40589 257897
rect 40623 257869 40651 257897
rect 40437 257807 40465 257835
rect 40499 257807 40527 257835
rect 40561 257807 40589 257835
rect 40623 257807 40651 257835
rect 40437 257745 40465 257773
rect 40499 257745 40527 257773
rect 40561 257745 40589 257773
rect 40623 257745 40651 257773
rect 47577 299162 47605 299190
rect 47639 299162 47667 299190
rect 47701 299162 47729 299190
rect 47763 299162 47791 299190
rect 47577 299100 47605 299128
rect 47639 299100 47667 299128
rect 47701 299100 47729 299128
rect 47763 299100 47791 299128
rect 47577 299038 47605 299066
rect 47639 299038 47667 299066
rect 47701 299038 47729 299066
rect 47763 299038 47791 299066
rect 47577 298976 47605 299004
rect 47639 298976 47667 299004
rect 47701 298976 47729 299004
rect 47763 298976 47791 299004
rect 47577 290931 47605 290959
rect 47639 290931 47667 290959
rect 47701 290931 47729 290959
rect 47763 290931 47791 290959
rect 47577 290869 47605 290897
rect 47639 290869 47667 290897
rect 47701 290869 47729 290897
rect 47763 290869 47791 290897
rect 47577 290807 47605 290835
rect 47639 290807 47667 290835
rect 47701 290807 47729 290835
rect 47763 290807 47791 290835
rect 47577 290745 47605 290773
rect 47639 290745 47667 290773
rect 47701 290745 47729 290773
rect 47763 290745 47791 290773
rect 47577 281931 47605 281959
rect 47639 281931 47667 281959
rect 47701 281931 47729 281959
rect 47763 281931 47791 281959
rect 47577 281869 47605 281897
rect 47639 281869 47667 281897
rect 47701 281869 47729 281897
rect 47763 281869 47791 281897
rect 47577 281807 47605 281835
rect 47639 281807 47667 281835
rect 47701 281807 47729 281835
rect 47763 281807 47791 281835
rect 47577 281745 47605 281773
rect 47639 281745 47667 281773
rect 47701 281745 47729 281773
rect 47763 281745 47791 281773
rect 47577 272931 47605 272959
rect 47639 272931 47667 272959
rect 47701 272931 47729 272959
rect 47763 272931 47791 272959
rect 47577 272869 47605 272897
rect 47639 272869 47667 272897
rect 47701 272869 47729 272897
rect 47763 272869 47791 272897
rect 47577 272807 47605 272835
rect 47639 272807 47667 272835
rect 47701 272807 47729 272835
rect 47763 272807 47791 272835
rect 47577 272745 47605 272773
rect 47639 272745 47667 272773
rect 47701 272745 47729 272773
rect 47763 272745 47791 272773
rect 47577 263931 47605 263959
rect 47639 263931 47667 263959
rect 47701 263931 47729 263959
rect 47763 263931 47791 263959
rect 47577 263869 47605 263897
rect 47639 263869 47667 263897
rect 47701 263869 47729 263897
rect 47763 263869 47791 263897
rect 47577 263807 47605 263835
rect 47639 263807 47667 263835
rect 47701 263807 47729 263835
rect 47763 263807 47791 263835
rect 47577 263745 47605 263773
rect 47639 263745 47667 263773
rect 47701 263745 47729 263773
rect 47763 263745 47791 263773
rect 47577 254931 47605 254959
rect 47639 254931 47667 254959
rect 47701 254931 47729 254959
rect 47763 254931 47791 254959
rect 47577 254869 47605 254897
rect 47639 254869 47667 254897
rect 47701 254869 47729 254897
rect 47763 254869 47791 254897
rect 47577 254807 47605 254835
rect 47639 254807 47667 254835
rect 47701 254807 47729 254835
rect 47763 254807 47791 254835
rect 47577 254745 47605 254773
rect 47639 254745 47667 254773
rect 47701 254745 47729 254773
rect 47763 254745 47791 254773
rect 49437 299642 49465 299670
rect 49499 299642 49527 299670
rect 49561 299642 49589 299670
rect 49623 299642 49651 299670
rect 49437 299580 49465 299608
rect 49499 299580 49527 299608
rect 49561 299580 49589 299608
rect 49623 299580 49651 299608
rect 49437 299518 49465 299546
rect 49499 299518 49527 299546
rect 49561 299518 49589 299546
rect 49623 299518 49651 299546
rect 49437 299456 49465 299484
rect 49499 299456 49527 299484
rect 49561 299456 49589 299484
rect 49623 299456 49651 299484
rect 49437 293931 49465 293959
rect 49499 293931 49527 293959
rect 49561 293931 49589 293959
rect 49623 293931 49651 293959
rect 49437 293869 49465 293897
rect 49499 293869 49527 293897
rect 49561 293869 49589 293897
rect 49623 293869 49651 293897
rect 49437 293807 49465 293835
rect 49499 293807 49527 293835
rect 49561 293807 49589 293835
rect 49623 293807 49651 293835
rect 49437 293745 49465 293773
rect 49499 293745 49527 293773
rect 49561 293745 49589 293773
rect 49623 293745 49651 293773
rect 49437 284931 49465 284959
rect 49499 284931 49527 284959
rect 49561 284931 49589 284959
rect 49623 284931 49651 284959
rect 49437 284869 49465 284897
rect 49499 284869 49527 284897
rect 49561 284869 49589 284897
rect 49623 284869 49651 284897
rect 49437 284807 49465 284835
rect 49499 284807 49527 284835
rect 49561 284807 49589 284835
rect 49623 284807 49651 284835
rect 49437 284745 49465 284773
rect 49499 284745 49527 284773
rect 49561 284745 49589 284773
rect 49623 284745 49651 284773
rect 49437 275931 49465 275959
rect 49499 275931 49527 275959
rect 49561 275931 49589 275959
rect 49623 275931 49651 275959
rect 49437 275869 49465 275897
rect 49499 275869 49527 275897
rect 49561 275869 49589 275897
rect 49623 275869 49651 275897
rect 49437 275807 49465 275835
rect 49499 275807 49527 275835
rect 49561 275807 49589 275835
rect 49623 275807 49651 275835
rect 49437 275745 49465 275773
rect 49499 275745 49527 275773
rect 49561 275745 49589 275773
rect 49623 275745 49651 275773
rect 49437 266931 49465 266959
rect 49499 266931 49527 266959
rect 49561 266931 49589 266959
rect 49623 266931 49651 266959
rect 49437 266869 49465 266897
rect 49499 266869 49527 266897
rect 49561 266869 49589 266897
rect 49623 266869 49651 266897
rect 49437 266807 49465 266835
rect 49499 266807 49527 266835
rect 49561 266807 49589 266835
rect 49623 266807 49651 266835
rect 49437 266745 49465 266773
rect 49499 266745 49527 266773
rect 49561 266745 49589 266773
rect 49623 266745 49651 266773
rect 49437 257931 49465 257959
rect 49499 257931 49527 257959
rect 49561 257931 49589 257959
rect 49623 257931 49651 257959
rect 49437 257869 49465 257897
rect 49499 257869 49527 257897
rect 49561 257869 49589 257897
rect 49623 257869 49651 257897
rect 49437 257807 49465 257835
rect 49499 257807 49527 257835
rect 49561 257807 49589 257835
rect 49623 257807 49651 257835
rect 49437 257745 49465 257773
rect 49499 257745 49527 257773
rect 49561 257745 49589 257773
rect 49623 257745 49651 257773
rect 56577 299162 56605 299190
rect 56639 299162 56667 299190
rect 56701 299162 56729 299190
rect 56763 299162 56791 299190
rect 56577 299100 56605 299128
rect 56639 299100 56667 299128
rect 56701 299100 56729 299128
rect 56763 299100 56791 299128
rect 56577 299038 56605 299066
rect 56639 299038 56667 299066
rect 56701 299038 56729 299066
rect 56763 299038 56791 299066
rect 56577 298976 56605 299004
rect 56639 298976 56667 299004
rect 56701 298976 56729 299004
rect 56763 298976 56791 299004
rect 56577 290931 56605 290959
rect 56639 290931 56667 290959
rect 56701 290931 56729 290959
rect 56763 290931 56791 290959
rect 56577 290869 56605 290897
rect 56639 290869 56667 290897
rect 56701 290869 56729 290897
rect 56763 290869 56791 290897
rect 56577 290807 56605 290835
rect 56639 290807 56667 290835
rect 56701 290807 56729 290835
rect 56763 290807 56791 290835
rect 56577 290745 56605 290773
rect 56639 290745 56667 290773
rect 56701 290745 56729 290773
rect 56763 290745 56791 290773
rect 56577 281931 56605 281959
rect 56639 281931 56667 281959
rect 56701 281931 56729 281959
rect 56763 281931 56791 281959
rect 56577 281869 56605 281897
rect 56639 281869 56667 281897
rect 56701 281869 56729 281897
rect 56763 281869 56791 281897
rect 56577 281807 56605 281835
rect 56639 281807 56667 281835
rect 56701 281807 56729 281835
rect 56763 281807 56791 281835
rect 56577 281745 56605 281773
rect 56639 281745 56667 281773
rect 56701 281745 56729 281773
rect 56763 281745 56791 281773
rect 56577 272931 56605 272959
rect 56639 272931 56667 272959
rect 56701 272931 56729 272959
rect 56763 272931 56791 272959
rect 56577 272869 56605 272897
rect 56639 272869 56667 272897
rect 56701 272869 56729 272897
rect 56763 272869 56791 272897
rect 56577 272807 56605 272835
rect 56639 272807 56667 272835
rect 56701 272807 56729 272835
rect 56763 272807 56791 272835
rect 56577 272745 56605 272773
rect 56639 272745 56667 272773
rect 56701 272745 56729 272773
rect 56763 272745 56791 272773
rect 56577 263931 56605 263959
rect 56639 263931 56667 263959
rect 56701 263931 56729 263959
rect 56763 263931 56791 263959
rect 56577 263869 56605 263897
rect 56639 263869 56667 263897
rect 56701 263869 56729 263897
rect 56763 263869 56791 263897
rect 56577 263807 56605 263835
rect 56639 263807 56667 263835
rect 56701 263807 56729 263835
rect 56763 263807 56791 263835
rect 56577 263745 56605 263773
rect 56639 263745 56667 263773
rect 56701 263745 56729 263773
rect 56763 263745 56791 263773
rect 56577 254931 56605 254959
rect 56639 254931 56667 254959
rect 56701 254931 56729 254959
rect 56763 254931 56791 254959
rect 56577 254869 56605 254897
rect 56639 254869 56667 254897
rect 56701 254869 56729 254897
rect 56763 254869 56791 254897
rect 56577 254807 56605 254835
rect 56639 254807 56667 254835
rect 56701 254807 56729 254835
rect 56763 254807 56791 254835
rect 56577 254745 56605 254773
rect 56639 254745 56667 254773
rect 56701 254745 56729 254773
rect 56763 254745 56791 254773
rect 58437 299642 58465 299670
rect 58499 299642 58527 299670
rect 58561 299642 58589 299670
rect 58623 299642 58651 299670
rect 58437 299580 58465 299608
rect 58499 299580 58527 299608
rect 58561 299580 58589 299608
rect 58623 299580 58651 299608
rect 58437 299518 58465 299546
rect 58499 299518 58527 299546
rect 58561 299518 58589 299546
rect 58623 299518 58651 299546
rect 58437 299456 58465 299484
rect 58499 299456 58527 299484
rect 58561 299456 58589 299484
rect 58623 299456 58651 299484
rect 58437 293931 58465 293959
rect 58499 293931 58527 293959
rect 58561 293931 58589 293959
rect 58623 293931 58651 293959
rect 58437 293869 58465 293897
rect 58499 293869 58527 293897
rect 58561 293869 58589 293897
rect 58623 293869 58651 293897
rect 58437 293807 58465 293835
rect 58499 293807 58527 293835
rect 58561 293807 58589 293835
rect 58623 293807 58651 293835
rect 58437 293745 58465 293773
rect 58499 293745 58527 293773
rect 58561 293745 58589 293773
rect 58623 293745 58651 293773
rect 58437 284931 58465 284959
rect 58499 284931 58527 284959
rect 58561 284931 58589 284959
rect 58623 284931 58651 284959
rect 58437 284869 58465 284897
rect 58499 284869 58527 284897
rect 58561 284869 58589 284897
rect 58623 284869 58651 284897
rect 58437 284807 58465 284835
rect 58499 284807 58527 284835
rect 58561 284807 58589 284835
rect 58623 284807 58651 284835
rect 58437 284745 58465 284773
rect 58499 284745 58527 284773
rect 58561 284745 58589 284773
rect 58623 284745 58651 284773
rect 58437 275931 58465 275959
rect 58499 275931 58527 275959
rect 58561 275931 58589 275959
rect 58623 275931 58651 275959
rect 58437 275869 58465 275897
rect 58499 275869 58527 275897
rect 58561 275869 58589 275897
rect 58623 275869 58651 275897
rect 58437 275807 58465 275835
rect 58499 275807 58527 275835
rect 58561 275807 58589 275835
rect 58623 275807 58651 275835
rect 58437 275745 58465 275773
rect 58499 275745 58527 275773
rect 58561 275745 58589 275773
rect 58623 275745 58651 275773
rect 58437 266931 58465 266959
rect 58499 266931 58527 266959
rect 58561 266931 58589 266959
rect 58623 266931 58651 266959
rect 58437 266869 58465 266897
rect 58499 266869 58527 266897
rect 58561 266869 58589 266897
rect 58623 266869 58651 266897
rect 58437 266807 58465 266835
rect 58499 266807 58527 266835
rect 58561 266807 58589 266835
rect 58623 266807 58651 266835
rect 58437 266745 58465 266773
rect 58499 266745 58527 266773
rect 58561 266745 58589 266773
rect 58623 266745 58651 266773
rect 58437 257931 58465 257959
rect 58499 257931 58527 257959
rect 58561 257931 58589 257959
rect 58623 257931 58651 257959
rect 58437 257869 58465 257897
rect 58499 257869 58527 257897
rect 58561 257869 58589 257897
rect 58623 257869 58651 257897
rect 58437 257807 58465 257835
rect 58499 257807 58527 257835
rect 58561 257807 58589 257835
rect 58623 257807 58651 257835
rect 58437 257745 58465 257773
rect 58499 257745 58527 257773
rect 58561 257745 58589 257773
rect 58623 257745 58651 257773
rect 65577 299162 65605 299190
rect 65639 299162 65667 299190
rect 65701 299162 65729 299190
rect 65763 299162 65791 299190
rect 65577 299100 65605 299128
rect 65639 299100 65667 299128
rect 65701 299100 65729 299128
rect 65763 299100 65791 299128
rect 65577 299038 65605 299066
rect 65639 299038 65667 299066
rect 65701 299038 65729 299066
rect 65763 299038 65791 299066
rect 65577 298976 65605 299004
rect 65639 298976 65667 299004
rect 65701 298976 65729 299004
rect 65763 298976 65791 299004
rect 65577 290931 65605 290959
rect 65639 290931 65667 290959
rect 65701 290931 65729 290959
rect 65763 290931 65791 290959
rect 65577 290869 65605 290897
rect 65639 290869 65667 290897
rect 65701 290869 65729 290897
rect 65763 290869 65791 290897
rect 65577 290807 65605 290835
rect 65639 290807 65667 290835
rect 65701 290807 65729 290835
rect 65763 290807 65791 290835
rect 65577 290745 65605 290773
rect 65639 290745 65667 290773
rect 65701 290745 65729 290773
rect 65763 290745 65791 290773
rect 65577 281931 65605 281959
rect 65639 281931 65667 281959
rect 65701 281931 65729 281959
rect 65763 281931 65791 281959
rect 65577 281869 65605 281897
rect 65639 281869 65667 281897
rect 65701 281869 65729 281897
rect 65763 281869 65791 281897
rect 65577 281807 65605 281835
rect 65639 281807 65667 281835
rect 65701 281807 65729 281835
rect 65763 281807 65791 281835
rect 65577 281745 65605 281773
rect 65639 281745 65667 281773
rect 65701 281745 65729 281773
rect 65763 281745 65791 281773
rect 65577 272931 65605 272959
rect 65639 272931 65667 272959
rect 65701 272931 65729 272959
rect 65763 272931 65791 272959
rect 65577 272869 65605 272897
rect 65639 272869 65667 272897
rect 65701 272869 65729 272897
rect 65763 272869 65791 272897
rect 65577 272807 65605 272835
rect 65639 272807 65667 272835
rect 65701 272807 65729 272835
rect 65763 272807 65791 272835
rect 65577 272745 65605 272773
rect 65639 272745 65667 272773
rect 65701 272745 65729 272773
rect 65763 272745 65791 272773
rect 65577 263931 65605 263959
rect 65639 263931 65667 263959
rect 65701 263931 65729 263959
rect 65763 263931 65791 263959
rect 65577 263869 65605 263897
rect 65639 263869 65667 263897
rect 65701 263869 65729 263897
rect 65763 263869 65791 263897
rect 65577 263807 65605 263835
rect 65639 263807 65667 263835
rect 65701 263807 65729 263835
rect 65763 263807 65791 263835
rect 65577 263745 65605 263773
rect 65639 263745 65667 263773
rect 65701 263745 65729 263773
rect 65763 263745 65791 263773
rect 65577 254931 65605 254959
rect 65639 254931 65667 254959
rect 65701 254931 65729 254959
rect 65763 254931 65791 254959
rect 65577 254869 65605 254897
rect 65639 254869 65667 254897
rect 65701 254869 65729 254897
rect 65763 254869 65791 254897
rect 65577 254807 65605 254835
rect 65639 254807 65667 254835
rect 65701 254807 65729 254835
rect 65763 254807 65791 254835
rect 65577 254745 65605 254773
rect 65639 254745 65667 254773
rect 65701 254745 65729 254773
rect 65763 254745 65791 254773
rect 67437 299642 67465 299670
rect 67499 299642 67527 299670
rect 67561 299642 67589 299670
rect 67623 299642 67651 299670
rect 67437 299580 67465 299608
rect 67499 299580 67527 299608
rect 67561 299580 67589 299608
rect 67623 299580 67651 299608
rect 67437 299518 67465 299546
rect 67499 299518 67527 299546
rect 67561 299518 67589 299546
rect 67623 299518 67651 299546
rect 67437 299456 67465 299484
rect 67499 299456 67527 299484
rect 67561 299456 67589 299484
rect 67623 299456 67651 299484
rect 67437 293931 67465 293959
rect 67499 293931 67527 293959
rect 67561 293931 67589 293959
rect 67623 293931 67651 293959
rect 67437 293869 67465 293897
rect 67499 293869 67527 293897
rect 67561 293869 67589 293897
rect 67623 293869 67651 293897
rect 67437 293807 67465 293835
rect 67499 293807 67527 293835
rect 67561 293807 67589 293835
rect 67623 293807 67651 293835
rect 67437 293745 67465 293773
rect 67499 293745 67527 293773
rect 67561 293745 67589 293773
rect 67623 293745 67651 293773
rect 67437 284931 67465 284959
rect 67499 284931 67527 284959
rect 67561 284931 67589 284959
rect 67623 284931 67651 284959
rect 67437 284869 67465 284897
rect 67499 284869 67527 284897
rect 67561 284869 67589 284897
rect 67623 284869 67651 284897
rect 67437 284807 67465 284835
rect 67499 284807 67527 284835
rect 67561 284807 67589 284835
rect 67623 284807 67651 284835
rect 67437 284745 67465 284773
rect 67499 284745 67527 284773
rect 67561 284745 67589 284773
rect 67623 284745 67651 284773
rect 67437 275931 67465 275959
rect 67499 275931 67527 275959
rect 67561 275931 67589 275959
rect 67623 275931 67651 275959
rect 67437 275869 67465 275897
rect 67499 275869 67527 275897
rect 67561 275869 67589 275897
rect 67623 275869 67651 275897
rect 67437 275807 67465 275835
rect 67499 275807 67527 275835
rect 67561 275807 67589 275835
rect 67623 275807 67651 275835
rect 67437 275745 67465 275773
rect 67499 275745 67527 275773
rect 67561 275745 67589 275773
rect 67623 275745 67651 275773
rect 67437 266931 67465 266959
rect 67499 266931 67527 266959
rect 67561 266931 67589 266959
rect 67623 266931 67651 266959
rect 67437 266869 67465 266897
rect 67499 266869 67527 266897
rect 67561 266869 67589 266897
rect 67623 266869 67651 266897
rect 67437 266807 67465 266835
rect 67499 266807 67527 266835
rect 67561 266807 67589 266835
rect 67623 266807 67651 266835
rect 67437 266745 67465 266773
rect 67499 266745 67527 266773
rect 67561 266745 67589 266773
rect 67623 266745 67651 266773
rect 67437 257931 67465 257959
rect 67499 257931 67527 257959
rect 67561 257931 67589 257959
rect 67623 257931 67651 257959
rect 67437 257869 67465 257897
rect 67499 257869 67527 257897
rect 67561 257869 67589 257897
rect 67623 257869 67651 257897
rect 67437 257807 67465 257835
rect 67499 257807 67527 257835
rect 67561 257807 67589 257835
rect 67623 257807 67651 257835
rect 67437 257745 67465 257773
rect 67499 257745 67527 257773
rect 67561 257745 67589 257773
rect 67623 257745 67651 257773
rect 74577 299162 74605 299190
rect 74639 299162 74667 299190
rect 74701 299162 74729 299190
rect 74763 299162 74791 299190
rect 74577 299100 74605 299128
rect 74639 299100 74667 299128
rect 74701 299100 74729 299128
rect 74763 299100 74791 299128
rect 74577 299038 74605 299066
rect 74639 299038 74667 299066
rect 74701 299038 74729 299066
rect 74763 299038 74791 299066
rect 74577 298976 74605 299004
rect 74639 298976 74667 299004
rect 74701 298976 74729 299004
rect 74763 298976 74791 299004
rect 74577 290931 74605 290959
rect 74639 290931 74667 290959
rect 74701 290931 74729 290959
rect 74763 290931 74791 290959
rect 74577 290869 74605 290897
rect 74639 290869 74667 290897
rect 74701 290869 74729 290897
rect 74763 290869 74791 290897
rect 74577 290807 74605 290835
rect 74639 290807 74667 290835
rect 74701 290807 74729 290835
rect 74763 290807 74791 290835
rect 74577 290745 74605 290773
rect 74639 290745 74667 290773
rect 74701 290745 74729 290773
rect 74763 290745 74791 290773
rect 74577 281931 74605 281959
rect 74639 281931 74667 281959
rect 74701 281931 74729 281959
rect 74763 281931 74791 281959
rect 74577 281869 74605 281897
rect 74639 281869 74667 281897
rect 74701 281869 74729 281897
rect 74763 281869 74791 281897
rect 74577 281807 74605 281835
rect 74639 281807 74667 281835
rect 74701 281807 74729 281835
rect 74763 281807 74791 281835
rect 74577 281745 74605 281773
rect 74639 281745 74667 281773
rect 74701 281745 74729 281773
rect 74763 281745 74791 281773
rect 74577 272931 74605 272959
rect 74639 272931 74667 272959
rect 74701 272931 74729 272959
rect 74763 272931 74791 272959
rect 74577 272869 74605 272897
rect 74639 272869 74667 272897
rect 74701 272869 74729 272897
rect 74763 272869 74791 272897
rect 74577 272807 74605 272835
rect 74639 272807 74667 272835
rect 74701 272807 74729 272835
rect 74763 272807 74791 272835
rect 74577 272745 74605 272773
rect 74639 272745 74667 272773
rect 74701 272745 74729 272773
rect 74763 272745 74791 272773
rect 74577 263931 74605 263959
rect 74639 263931 74667 263959
rect 74701 263931 74729 263959
rect 74763 263931 74791 263959
rect 74577 263869 74605 263897
rect 74639 263869 74667 263897
rect 74701 263869 74729 263897
rect 74763 263869 74791 263897
rect 74577 263807 74605 263835
rect 74639 263807 74667 263835
rect 74701 263807 74729 263835
rect 74763 263807 74791 263835
rect 74577 263745 74605 263773
rect 74639 263745 74667 263773
rect 74701 263745 74729 263773
rect 74763 263745 74791 263773
rect 74577 254931 74605 254959
rect 74639 254931 74667 254959
rect 74701 254931 74729 254959
rect 74763 254931 74791 254959
rect 74577 254869 74605 254897
rect 74639 254869 74667 254897
rect 74701 254869 74729 254897
rect 74763 254869 74791 254897
rect 74577 254807 74605 254835
rect 74639 254807 74667 254835
rect 74701 254807 74729 254835
rect 74763 254807 74791 254835
rect 74577 254745 74605 254773
rect 74639 254745 74667 254773
rect 74701 254745 74729 254773
rect 74763 254745 74791 254773
rect 76437 299642 76465 299670
rect 76499 299642 76527 299670
rect 76561 299642 76589 299670
rect 76623 299642 76651 299670
rect 76437 299580 76465 299608
rect 76499 299580 76527 299608
rect 76561 299580 76589 299608
rect 76623 299580 76651 299608
rect 76437 299518 76465 299546
rect 76499 299518 76527 299546
rect 76561 299518 76589 299546
rect 76623 299518 76651 299546
rect 76437 299456 76465 299484
rect 76499 299456 76527 299484
rect 76561 299456 76589 299484
rect 76623 299456 76651 299484
rect 76437 293931 76465 293959
rect 76499 293931 76527 293959
rect 76561 293931 76589 293959
rect 76623 293931 76651 293959
rect 76437 293869 76465 293897
rect 76499 293869 76527 293897
rect 76561 293869 76589 293897
rect 76623 293869 76651 293897
rect 76437 293807 76465 293835
rect 76499 293807 76527 293835
rect 76561 293807 76589 293835
rect 76623 293807 76651 293835
rect 76437 293745 76465 293773
rect 76499 293745 76527 293773
rect 76561 293745 76589 293773
rect 76623 293745 76651 293773
rect 76437 284931 76465 284959
rect 76499 284931 76527 284959
rect 76561 284931 76589 284959
rect 76623 284931 76651 284959
rect 76437 284869 76465 284897
rect 76499 284869 76527 284897
rect 76561 284869 76589 284897
rect 76623 284869 76651 284897
rect 76437 284807 76465 284835
rect 76499 284807 76527 284835
rect 76561 284807 76589 284835
rect 76623 284807 76651 284835
rect 76437 284745 76465 284773
rect 76499 284745 76527 284773
rect 76561 284745 76589 284773
rect 76623 284745 76651 284773
rect 76437 275931 76465 275959
rect 76499 275931 76527 275959
rect 76561 275931 76589 275959
rect 76623 275931 76651 275959
rect 76437 275869 76465 275897
rect 76499 275869 76527 275897
rect 76561 275869 76589 275897
rect 76623 275869 76651 275897
rect 76437 275807 76465 275835
rect 76499 275807 76527 275835
rect 76561 275807 76589 275835
rect 76623 275807 76651 275835
rect 76437 275745 76465 275773
rect 76499 275745 76527 275773
rect 76561 275745 76589 275773
rect 76623 275745 76651 275773
rect 76437 266931 76465 266959
rect 76499 266931 76527 266959
rect 76561 266931 76589 266959
rect 76623 266931 76651 266959
rect 76437 266869 76465 266897
rect 76499 266869 76527 266897
rect 76561 266869 76589 266897
rect 76623 266869 76651 266897
rect 76437 266807 76465 266835
rect 76499 266807 76527 266835
rect 76561 266807 76589 266835
rect 76623 266807 76651 266835
rect 76437 266745 76465 266773
rect 76499 266745 76527 266773
rect 76561 266745 76589 266773
rect 76623 266745 76651 266773
rect 76437 257931 76465 257959
rect 76499 257931 76527 257959
rect 76561 257931 76589 257959
rect 76623 257931 76651 257959
rect 76437 257869 76465 257897
rect 76499 257869 76527 257897
rect 76561 257869 76589 257897
rect 76623 257869 76651 257897
rect 76437 257807 76465 257835
rect 76499 257807 76527 257835
rect 76561 257807 76589 257835
rect 76623 257807 76651 257835
rect 76437 257745 76465 257773
rect 76499 257745 76527 257773
rect 76561 257745 76589 257773
rect 76623 257745 76651 257773
rect 83577 299162 83605 299190
rect 83639 299162 83667 299190
rect 83701 299162 83729 299190
rect 83763 299162 83791 299190
rect 83577 299100 83605 299128
rect 83639 299100 83667 299128
rect 83701 299100 83729 299128
rect 83763 299100 83791 299128
rect 83577 299038 83605 299066
rect 83639 299038 83667 299066
rect 83701 299038 83729 299066
rect 83763 299038 83791 299066
rect 83577 298976 83605 299004
rect 83639 298976 83667 299004
rect 83701 298976 83729 299004
rect 83763 298976 83791 299004
rect 83577 290931 83605 290959
rect 83639 290931 83667 290959
rect 83701 290931 83729 290959
rect 83763 290931 83791 290959
rect 83577 290869 83605 290897
rect 83639 290869 83667 290897
rect 83701 290869 83729 290897
rect 83763 290869 83791 290897
rect 83577 290807 83605 290835
rect 83639 290807 83667 290835
rect 83701 290807 83729 290835
rect 83763 290807 83791 290835
rect 83577 290745 83605 290773
rect 83639 290745 83667 290773
rect 83701 290745 83729 290773
rect 83763 290745 83791 290773
rect 83577 281931 83605 281959
rect 83639 281931 83667 281959
rect 83701 281931 83729 281959
rect 83763 281931 83791 281959
rect 83577 281869 83605 281897
rect 83639 281869 83667 281897
rect 83701 281869 83729 281897
rect 83763 281869 83791 281897
rect 83577 281807 83605 281835
rect 83639 281807 83667 281835
rect 83701 281807 83729 281835
rect 83763 281807 83791 281835
rect 83577 281745 83605 281773
rect 83639 281745 83667 281773
rect 83701 281745 83729 281773
rect 83763 281745 83791 281773
rect 83577 272931 83605 272959
rect 83639 272931 83667 272959
rect 83701 272931 83729 272959
rect 83763 272931 83791 272959
rect 83577 272869 83605 272897
rect 83639 272869 83667 272897
rect 83701 272869 83729 272897
rect 83763 272869 83791 272897
rect 83577 272807 83605 272835
rect 83639 272807 83667 272835
rect 83701 272807 83729 272835
rect 83763 272807 83791 272835
rect 83577 272745 83605 272773
rect 83639 272745 83667 272773
rect 83701 272745 83729 272773
rect 83763 272745 83791 272773
rect 83577 263931 83605 263959
rect 83639 263931 83667 263959
rect 83701 263931 83729 263959
rect 83763 263931 83791 263959
rect 83577 263869 83605 263897
rect 83639 263869 83667 263897
rect 83701 263869 83729 263897
rect 83763 263869 83791 263897
rect 83577 263807 83605 263835
rect 83639 263807 83667 263835
rect 83701 263807 83729 263835
rect 83763 263807 83791 263835
rect 83577 263745 83605 263773
rect 83639 263745 83667 263773
rect 83701 263745 83729 263773
rect 83763 263745 83791 263773
rect 83577 254931 83605 254959
rect 83639 254931 83667 254959
rect 83701 254931 83729 254959
rect 83763 254931 83791 254959
rect 83577 254869 83605 254897
rect 83639 254869 83667 254897
rect 83701 254869 83729 254897
rect 83763 254869 83791 254897
rect 83577 254807 83605 254835
rect 83639 254807 83667 254835
rect 83701 254807 83729 254835
rect 83763 254807 83791 254835
rect 83577 254745 83605 254773
rect 83639 254745 83667 254773
rect 83701 254745 83729 254773
rect 83763 254745 83791 254773
rect 85437 299642 85465 299670
rect 85499 299642 85527 299670
rect 85561 299642 85589 299670
rect 85623 299642 85651 299670
rect 85437 299580 85465 299608
rect 85499 299580 85527 299608
rect 85561 299580 85589 299608
rect 85623 299580 85651 299608
rect 85437 299518 85465 299546
rect 85499 299518 85527 299546
rect 85561 299518 85589 299546
rect 85623 299518 85651 299546
rect 85437 299456 85465 299484
rect 85499 299456 85527 299484
rect 85561 299456 85589 299484
rect 85623 299456 85651 299484
rect 85437 293931 85465 293959
rect 85499 293931 85527 293959
rect 85561 293931 85589 293959
rect 85623 293931 85651 293959
rect 85437 293869 85465 293897
rect 85499 293869 85527 293897
rect 85561 293869 85589 293897
rect 85623 293869 85651 293897
rect 85437 293807 85465 293835
rect 85499 293807 85527 293835
rect 85561 293807 85589 293835
rect 85623 293807 85651 293835
rect 85437 293745 85465 293773
rect 85499 293745 85527 293773
rect 85561 293745 85589 293773
rect 85623 293745 85651 293773
rect 85437 284931 85465 284959
rect 85499 284931 85527 284959
rect 85561 284931 85589 284959
rect 85623 284931 85651 284959
rect 85437 284869 85465 284897
rect 85499 284869 85527 284897
rect 85561 284869 85589 284897
rect 85623 284869 85651 284897
rect 85437 284807 85465 284835
rect 85499 284807 85527 284835
rect 85561 284807 85589 284835
rect 85623 284807 85651 284835
rect 85437 284745 85465 284773
rect 85499 284745 85527 284773
rect 85561 284745 85589 284773
rect 85623 284745 85651 284773
rect 85437 275931 85465 275959
rect 85499 275931 85527 275959
rect 85561 275931 85589 275959
rect 85623 275931 85651 275959
rect 85437 275869 85465 275897
rect 85499 275869 85527 275897
rect 85561 275869 85589 275897
rect 85623 275869 85651 275897
rect 85437 275807 85465 275835
rect 85499 275807 85527 275835
rect 85561 275807 85589 275835
rect 85623 275807 85651 275835
rect 85437 275745 85465 275773
rect 85499 275745 85527 275773
rect 85561 275745 85589 275773
rect 85623 275745 85651 275773
rect 85437 266931 85465 266959
rect 85499 266931 85527 266959
rect 85561 266931 85589 266959
rect 85623 266931 85651 266959
rect 85437 266869 85465 266897
rect 85499 266869 85527 266897
rect 85561 266869 85589 266897
rect 85623 266869 85651 266897
rect 85437 266807 85465 266835
rect 85499 266807 85527 266835
rect 85561 266807 85589 266835
rect 85623 266807 85651 266835
rect 85437 266745 85465 266773
rect 85499 266745 85527 266773
rect 85561 266745 85589 266773
rect 85623 266745 85651 266773
rect 85437 257931 85465 257959
rect 85499 257931 85527 257959
rect 85561 257931 85589 257959
rect 85623 257931 85651 257959
rect 85437 257869 85465 257897
rect 85499 257869 85527 257897
rect 85561 257869 85589 257897
rect 85623 257869 85651 257897
rect 85437 257807 85465 257835
rect 85499 257807 85527 257835
rect 85561 257807 85589 257835
rect 85623 257807 85651 257835
rect 85437 257745 85465 257773
rect 85499 257745 85527 257773
rect 85561 257745 85589 257773
rect 85623 257745 85651 257773
rect 92577 299162 92605 299190
rect 92639 299162 92667 299190
rect 92701 299162 92729 299190
rect 92763 299162 92791 299190
rect 92577 299100 92605 299128
rect 92639 299100 92667 299128
rect 92701 299100 92729 299128
rect 92763 299100 92791 299128
rect 92577 299038 92605 299066
rect 92639 299038 92667 299066
rect 92701 299038 92729 299066
rect 92763 299038 92791 299066
rect 92577 298976 92605 299004
rect 92639 298976 92667 299004
rect 92701 298976 92729 299004
rect 92763 298976 92791 299004
rect 92577 290931 92605 290959
rect 92639 290931 92667 290959
rect 92701 290931 92729 290959
rect 92763 290931 92791 290959
rect 92577 290869 92605 290897
rect 92639 290869 92667 290897
rect 92701 290869 92729 290897
rect 92763 290869 92791 290897
rect 92577 290807 92605 290835
rect 92639 290807 92667 290835
rect 92701 290807 92729 290835
rect 92763 290807 92791 290835
rect 92577 290745 92605 290773
rect 92639 290745 92667 290773
rect 92701 290745 92729 290773
rect 92763 290745 92791 290773
rect 92577 281931 92605 281959
rect 92639 281931 92667 281959
rect 92701 281931 92729 281959
rect 92763 281931 92791 281959
rect 92577 281869 92605 281897
rect 92639 281869 92667 281897
rect 92701 281869 92729 281897
rect 92763 281869 92791 281897
rect 92577 281807 92605 281835
rect 92639 281807 92667 281835
rect 92701 281807 92729 281835
rect 92763 281807 92791 281835
rect 92577 281745 92605 281773
rect 92639 281745 92667 281773
rect 92701 281745 92729 281773
rect 92763 281745 92791 281773
rect 92577 272931 92605 272959
rect 92639 272931 92667 272959
rect 92701 272931 92729 272959
rect 92763 272931 92791 272959
rect 92577 272869 92605 272897
rect 92639 272869 92667 272897
rect 92701 272869 92729 272897
rect 92763 272869 92791 272897
rect 92577 272807 92605 272835
rect 92639 272807 92667 272835
rect 92701 272807 92729 272835
rect 92763 272807 92791 272835
rect 92577 272745 92605 272773
rect 92639 272745 92667 272773
rect 92701 272745 92729 272773
rect 92763 272745 92791 272773
rect 92577 263931 92605 263959
rect 92639 263931 92667 263959
rect 92701 263931 92729 263959
rect 92763 263931 92791 263959
rect 92577 263869 92605 263897
rect 92639 263869 92667 263897
rect 92701 263869 92729 263897
rect 92763 263869 92791 263897
rect 92577 263807 92605 263835
rect 92639 263807 92667 263835
rect 92701 263807 92729 263835
rect 92763 263807 92791 263835
rect 92577 263745 92605 263773
rect 92639 263745 92667 263773
rect 92701 263745 92729 263773
rect 92763 263745 92791 263773
rect 92577 254931 92605 254959
rect 92639 254931 92667 254959
rect 92701 254931 92729 254959
rect 92763 254931 92791 254959
rect 92577 254869 92605 254897
rect 92639 254869 92667 254897
rect 92701 254869 92729 254897
rect 92763 254869 92791 254897
rect 92577 254807 92605 254835
rect 92639 254807 92667 254835
rect 92701 254807 92729 254835
rect 92763 254807 92791 254835
rect 92577 254745 92605 254773
rect 92639 254745 92667 254773
rect 92701 254745 92729 254773
rect 92763 254745 92791 254773
rect 94437 299642 94465 299670
rect 94499 299642 94527 299670
rect 94561 299642 94589 299670
rect 94623 299642 94651 299670
rect 94437 299580 94465 299608
rect 94499 299580 94527 299608
rect 94561 299580 94589 299608
rect 94623 299580 94651 299608
rect 94437 299518 94465 299546
rect 94499 299518 94527 299546
rect 94561 299518 94589 299546
rect 94623 299518 94651 299546
rect 94437 299456 94465 299484
rect 94499 299456 94527 299484
rect 94561 299456 94589 299484
rect 94623 299456 94651 299484
rect 94437 293931 94465 293959
rect 94499 293931 94527 293959
rect 94561 293931 94589 293959
rect 94623 293931 94651 293959
rect 94437 293869 94465 293897
rect 94499 293869 94527 293897
rect 94561 293869 94589 293897
rect 94623 293869 94651 293897
rect 94437 293807 94465 293835
rect 94499 293807 94527 293835
rect 94561 293807 94589 293835
rect 94623 293807 94651 293835
rect 94437 293745 94465 293773
rect 94499 293745 94527 293773
rect 94561 293745 94589 293773
rect 94623 293745 94651 293773
rect 94437 284931 94465 284959
rect 94499 284931 94527 284959
rect 94561 284931 94589 284959
rect 94623 284931 94651 284959
rect 94437 284869 94465 284897
rect 94499 284869 94527 284897
rect 94561 284869 94589 284897
rect 94623 284869 94651 284897
rect 94437 284807 94465 284835
rect 94499 284807 94527 284835
rect 94561 284807 94589 284835
rect 94623 284807 94651 284835
rect 94437 284745 94465 284773
rect 94499 284745 94527 284773
rect 94561 284745 94589 284773
rect 94623 284745 94651 284773
rect 94437 275931 94465 275959
rect 94499 275931 94527 275959
rect 94561 275931 94589 275959
rect 94623 275931 94651 275959
rect 94437 275869 94465 275897
rect 94499 275869 94527 275897
rect 94561 275869 94589 275897
rect 94623 275869 94651 275897
rect 94437 275807 94465 275835
rect 94499 275807 94527 275835
rect 94561 275807 94589 275835
rect 94623 275807 94651 275835
rect 94437 275745 94465 275773
rect 94499 275745 94527 275773
rect 94561 275745 94589 275773
rect 94623 275745 94651 275773
rect 94437 266931 94465 266959
rect 94499 266931 94527 266959
rect 94561 266931 94589 266959
rect 94623 266931 94651 266959
rect 94437 266869 94465 266897
rect 94499 266869 94527 266897
rect 94561 266869 94589 266897
rect 94623 266869 94651 266897
rect 94437 266807 94465 266835
rect 94499 266807 94527 266835
rect 94561 266807 94589 266835
rect 94623 266807 94651 266835
rect 94437 266745 94465 266773
rect 94499 266745 94527 266773
rect 94561 266745 94589 266773
rect 94623 266745 94651 266773
rect 94437 257931 94465 257959
rect 94499 257931 94527 257959
rect 94561 257931 94589 257959
rect 94623 257931 94651 257959
rect 94437 257869 94465 257897
rect 94499 257869 94527 257897
rect 94561 257869 94589 257897
rect 94623 257869 94651 257897
rect 94437 257807 94465 257835
rect 94499 257807 94527 257835
rect 94561 257807 94589 257835
rect 94623 257807 94651 257835
rect 94437 257745 94465 257773
rect 94499 257745 94527 257773
rect 94561 257745 94589 257773
rect 94623 257745 94651 257773
rect 101577 299162 101605 299190
rect 101639 299162 101667 299190
rect 101701 299162 101729 299190
rect 101763 299162 101791 299190
rect 101577 299100 101605 299128
rect 101639 299100 101667 299128
rect 101701 299100 101729 299128
rect 101763 299100 101791 299128
rect 101577 299038 101605 299066
rect 101639 299038 101667 299066
rect 101701 299038 101729 299066
rect 101763 299038 101791 299066
rect 101577 298976 101605 299004
rect 101639 298976 101667 299004
rect 101701 298976 101729 299004
rect 101763 298976 101791 299004
rect 101577 290931 101605 290959
rect 101639 290931 101667 290959
rect 101701 290931 101729 290959
rect 101763 290931 101791 290959
rect 101577 290869 101605 290897
rect 101639 290869 101667 290897
rect 101701 290869 101729 290897
rect 101763 290869 101791 290897
rect 101577 290807 101605 290835
rect 101639 290807 101667 290835
rect 101701 290807 101729 290835
rect 101763 290807 101791 290835
rect 101577 290745 101605 290773
rect 101639 290745 101667 290773
rect 101701 290745 101729 290773
rect 101763 290745 101791 290773
rect 101577 281931 101605 281959
rect 101639 281931 101667 281959
rect 101701 281931 101729 281959
rect 101763 281931 101791 281959
rect 101577 281869 101605 281897
rect 101639 281869 101667 281897
rect 101701 281869 101729 281897
rect 101763 281869 101791 281897
rect 101577 281807 101605 281835
rect 101639 281807 101667 281835
rect 101701 281807 101729 281835
rect 101763 281807 101791 281835
rect 101577 281745 101605 281773
rect 101639 281745 101667 281773
rect 101701 281745 101729 281773
rect 101763 281745 101791 281773
rect 101577 272931 101605 272959
rect 101639 272931 101667 272959
rect 101701 272931 101729 272959
rect 101763 272931 101791 272959
rect 101577 272869 101605 272897
rect 101639 272869 101667 272897
rect 101701 272869 101729 272897
rect 101763 272869 101791 272897
rect 101577 272807 101605 272835
rect 101639 272807 101667 272835
rect 101701 272807 101729 272835
rect 101763 272807 101791 272835
rect 101577 272745 101605 272773
rect 101639 272745 101667 272773
rect 101701 272745 101729 272773
rect 101763 272745 101791 272773
rect 101577 263931 101605 263959
rect 101639 263931 101667 263959
rect 101701 263931 101729 263959
rect 101763 263931 101791 263959
rect 101577 263869 101605 263897
rect 101639 263869 101667 263897
rect 101701 263869 101729 263897
rect 101763 263869 101791 263897
rect 101577 263807 101605 263835
rect 101639 263807 101667 263835
rect 101701 263807 101729 263835
rect 101763 263807 101791 263835
rect 101577 263745 101605 263773
rect 101639 263745 101667 263773
rect 101701 263745 101729 263773
rect 101763 263745 101791 263773
rect 101577 254931 101605 254959
rect 101639 254931 101667 254959
rect 101701 254931 101729 254959
rect 101763 254931 101791 254959
rect 101577 254869 101605 254897
rect 101639 254869 101667 254897
rect 101701 254869 101729 254897
rect 101763 254869 101791 254897
rect 101577 254807 101605 254835
rect 101639 254807 101667 254835
rect 101701 254807 101729 254835
rect 101763 254807 101791 254835
rect 101577 254745 101605 254773
rect 101639 254745 101667 254773
rect 101701 254745 101729 254773
rect 101763 254745 101791 254773
rect 103437 299642 103465 299670
rect 103499 299642 103527 299670
rect 103561 299642 103589 299670
rect 103623 299642 103651 299670
rect 103437 299580 103465 299608
rect 103499 299580 103527 299608
rect 103561 299580 103589 299608
rect 103623 299580 103651 299608
rect 103437 299518 103465 299546
rect 103499 299518 103527 299546
rect 103561 299518 103589 299546
rect 103623 299518 103651 299546
rect 103437 299456 103465 299484
rect 103499 299456 103527 299484
rect 103561 299456 103589 299484
rect 103623 299456 103651 299484
rect 103437 293931 103465 293959
rect 103499 293931 103527 293959
rect 103561 293931 103589 293959
rect 103623 293931 103651 293959
rect 103437 293869 103465 293897
rect 103499 293869 103527 293897
rect 103561 293869 103589 293897
rect 103623 293869 103651 293897
rect 103437 293807 103465 293835
rect 103499 293807 103527 293835
rect 103561 293807 103589 293835
rect 103623 293807 103651 293835
rect 103437 293745 103465 293773
rect 103499 293745 103527 293773
rect 103561 293745 103589 293773
rect 103623 293745 103651 293773
rect 103437 284931 103465 284959
rect 103499 284931 103527 284959
rect 103561 284931 103589 284959
rect 103623 284931 103651 284959
rect 103437 284869 103465 284897
rect 103499 284869 103527 284897
rect 103561 284869 103589 284897
rect 103623 284869 103651 284897
rect 103437 284807 103465 284835
rect 103499 284807 103527 284835
rect 103561 284807 103589 284835
rect 103623 284807 103651 284835
rect 103437 284745 103465 284773
rect 103499 284745 103527 284773
rect 103561 284745 103589 284773
rect 103623 284745 103651 284773
rect 103437 275931 103465 275959
rect 103499 275931 103527 275959
rect 103561 275931 103589 275959
rect 103623 275931 103651 275959
rect 103437 275869 103465 275897
rect 103499 275869 103527 275897
rect 103561 275869 103589 275897
rect 103623 275869 103651 275897
rect 103437 275807 103465 275835
rect 103499 275807 103527 275835
rect 103561 275807 103589 275835
rect 103623 275807 103651 275835
rect 103437 275745 103465 275773
rect 103499 275745 103527 275773
rect 103561 275745 103589 275773
rect 103623 275745 103651 275773
rect 103437 266931 103465 266959
rect 103499 266931 103527 266959
rect 103561 266931 103589 266959
rect 103623 266931 103651 266959
rect 103437 266869 103465 266897
rect 103499 266869 103527 266897
rect 103561 266869 103589 266897
rect 103623 266869 103651 266897
rect 103437 266807 103465 266835
rect 103499 266807 103527 266835
rect 103561 266807 103589 266835
rect 103623 266807 103651 266835
rect 103437 266745 103465 266773
rect 103499 266745 103527 266773
rect 103561 266745 103589 266773
rect 103623 266745 103651 266773
rect 103437 257931 103465 257959
rect 103499 257931 103527 257959
rect 103561 257931 103589 257959
rect 103623 257931 103651 257959
rect 103437 257869 103465 257897
rect 103499 257869 103527 257897
rect 103561 257869 103589 257897
rect 103623 257869 103651 257897
rect 103437 257807 103465 257835
rect 103499 257807 103527 257835
rect 103561 257807 103589 257835
rect 103623 257807 103651 257835
rect 103437 257745 103465 257773
rect 103499 257745 103527 257773
rect 103561 257745 103589 257773
rect 103623 257745 103651 257773
rect 110577 299162 110605 299190
rect 110639 299162 110667 299190
rect 110701 299162 110729 299190
rect 110763 299162 110791 299190
rect 110577 299100 110605 299128
rect 110639 299100 110667 299128
rect 110701 299100 110729 299128
rect 110763 299100 110791 299128
rect 110577 299038 110605 299066
rect 110639 299038 110667 299066
rect 110701 299038 110729 299066
rect 110763 299038 110791 299066
rect 110577 298976 110605 299004
rect 110639 298976 110667 299004
rect 110701 298976 110729 299004
rect 110763 298976 110791 299004
rect 110577 290931 110605 290959
rect 110639 290931 110667 290959
rect 110701 290931 110729 290959
rect 110763 290931 110791 290959
rect 110577 290869 110605 290897
rect 110639 290869 110667 290897
rect 110701 290869 110729 290897
rect 110763 290869 110791 290897
rect 110577 290807 110605 290835
rect 110639 290807 110667 290835
rect 110701 290807 110729 290835
rect 110763 290807 110791 290835
rect 110577 290745 110605 290773
rect 110639 290745 110667 290773
rect 110701 290745 110729 290773
rect 110763 290745 110791 290773
rect 110577 281931 110605 281959
rect 110639 281931 110667 281959
rect 110701 281931 110729 281959
rect 110763 281931 110791 281959
rect 110577 281869 110605 281897
rect 110639 281869 110667 281897
rect 110701 281869 110729 281897
rect 110763 281869 110791 281897
rect 110577 281807 110605 281835
rect 110639 281807 110667 281835
rect 110701 281807 110729 281835
rect 110763 281807 110791 281835
rect 110577 281745 110605 281773
rect 110639 281745 110667 281773
rect 110701 281745 110729 281773
rect 110763 281745 110791 281773
rect 110577 272931 110605 272959
rect 110639 272931 110667 272959
rect 110701 272931 110729 272959
rect 110763 272931 110791 272959
rect 110577 272869 110605 272897
rect 110639 272869 110667 272897
rect 110701 272869 110729 272897
rect 110763 272869 110791 272897
rect 110577 272807 110605 272835
rect 110639 272807 110667 272835
rect 110701 272807 110729 272835
rect 110763 272807 110791 272835
rect 110577 272745 110605 272773
rect 110639 272745 110667 272773
rect 110701 272745 110729 272773
rect 110763 272745 110791 272773
rect 110577 263931 110605 263959
rect 110639 263931 110667 263959
rect 110701 263931 110729 263959
rect 110763 263931 110791 263959
rect 110577 263869 110605 263897
rect 110639 263869 110667 263897
rect 110701 263869 110729 263897
rect 110763 263869 110791 263897
rect 110577 263807 110605 263835
rect 110639 263807 110667 263835
rect 110701 263807 110729 263835
rect 110763 263807 110791 263835
rect 110577 263745 110605 263773
rect 110639 263745 110667 263773
rect 110701 263745 110729 263773
rect 110763 263745 110791 263773
rect 110577 254931 110605 254959
rect 110639 254931 110667 254959
rect 110701 254931 110729 254959
rect 110763 254931 110791 254959
rect 110577 254869 110605 254897
rect 110639 254869 110667 254897
rect 110701 254869 110729 254897
rect 110763 254869 110791 254897
rect 110577 254807 110605 254835
rect 110639 254807 110667 254835
rect 110701 254807 110729 254835
rect 110763 254807 110791 254835
rect 110577 254745 110605 254773
rect 110639 254745 110667 254773
rect 110701 254745 110729 254773
rect 110763 254745 110791 254773
rect 112437 299642 112465 299670
rect 112499 299642 112527 299670
rect 112561 299642 112589 299670
rect 112623 299642 112651 299670
rect 112437 299580 112465 299608
rect 112499 299580 112527 299608
rect 112561 299580 112589 299608
rect 112623 299580 112651 299608
rect 112437 299518 112465 299546
rect 112499 299518 112527 299546
rect 112561 299518 112589 299546
rect 112623 299518 112651 299546
rect 112437 299456 112465 299484
rect 112499 299456 112527 299484
rect 112561 299456 112589 299484
rect 112623 299456 112651 299484
rect 112437 293931 112465 293959
rect 112499 293931 112527 293959
rect 112561 293931 112589 293959
rect 112623 293931 112651 293959
rect 112437 293869 112465 293897
rect 112499 293869 112527 293897
rect 112561 293869 112589 293897
rect 112623 293869 112651 293897
rect 112437 293807 112465 293835
rect 112499 293807 112527 293835
rect 112561 293807 112589 293835
rect 112623 293807 112651 293835
rect 112437 293745 112465 293773
rect 112499 293745 112527 293773
rect 112561 293745 112589 293773
rect 112623 293745 112651 293773
rect 112437 284931 112465 284959
rect 112499 284931 112527 284959
rect 112561 284931 112589 284959
rect 112623 284931 112651 284959
rect 112437 284869 112465 284897
rect 112499 284869 112527 284897
rect 112561 284869 112589 284897
rect 112623 284869 112651 284897
rect 112437 284807 112465 284835
rect 112499 284807 112527 284835
rect 112561 284807 112589 284835
rect 112623 284807 112651 284835
rect 112437 284745 112465 284773
rect 112499 284745 112527 284773
rect 112561 284745 112589 284773
rect 112623 284745 112651 284773
rect 112437 275931 112465 275959
rect 112499 275931 112527 275959
rect 112561 275931 112589 275959
rect 112623 275931 112651 275959
rect 112437 275869 112465 275897
rect 112499 275869 112527 275897
rect 112561 275869 112589 275897
rect 112623 275869 112651 275897
rect 112437 275807 112465 275835
rect 112499 275807 112527 275835
rect 112561 275807 112589 275835
rect 112623 275807 112651 275835
rect 112437 275745 112465 275773
rect 112499 275745 112527 275773
rect 112561 275745 112589 275773
rect 112623 275745 112651 275773
rect 112437 266931 112465 266959
rect 112499 266931 112527 266959
rect 112561 266931 112589 266959
rect 112623 266931 112651 266959
rect 112437 266869 112465 266897
rect 112499 266869 112527 266897
rect 112561 266869 112589 266897
rect 112623 266869 112651 266897
rect 112437 266807 112465 266835
rect 112499 266807 112527 266835
rect 112561 266807 112589 266835
rect 112623 266807 112651 266835
rect 112437 266745 112465 266773
rect 112499 266745 112527 266773
rect 112561 266745 112589 266773
rect 112623 266745 112651 266773
rect 112437 257931 112465 257959
rect 112499 257931 112527 257959
rect 112561 257931 112589 257959
rect 112623 257931 112651 257959
rect 112437 257869 112465 257897
rect 112499 257869 112527 257897
rect 112561 257869 112589 257897
rect 112623 257869 112651 257897
rect 112437 257807 112465 257835
rect 112499 257807 112527 257835
rect 112561 257807 112589 257835
rect 112623 257807 112651 257835
rect 112437 257745 112465 257773
rect 112499 257745 112527 257773
rect 112561 257745 112589 257773
rect 112623 257745 112651 257773
rect 119577 299162 119605 299190
rect 119639 299162 119667 299190
rect 119701 299162 119729 299190
rect 119763 299162 119791 299190
rect 119577 299100 119605 299128
rect 119639 299100 119667 299128
rect 119701 299100 119729 299128
rect 119763 299100 119791 299128
rect 119577 299038 119605 299066
rect 119639 299038 119667 299066
rect 119701 299038 119729 299066
rect 119763 299038 119791 299066
rect 119577 298976 119605 299004
rect 119639 298976 119667 299004
rect 119701 298976 119729 299004
rect 119763 298976 119791 299004
rect 119577 290931 119605 290959
rect 119639 290931 119667 290959
rect 119701 290931 119729 290959
rect 119763 290931 119791 290959
rect 119577 290869 119605 290897
rect 119639 290869 119667 290897
rect 119701 290869 119729 290897
rect 119763 290869 119791 290897
rect 119577 290807 119605 290835
rect 119639 290807 119667 290835
rect 119701 290807 119729 290835
rect 119763 290807 119791 290835
rect 119577 290745 119605 290773
rect 119639 290745 119667 290773
rect 119701 290745 119729 290773
rect 119763 290745 119791 290773
rect 119577 281931 119605 281959
rect 119639 281931 119667 281959
rect 119701 281931 119729 281959
rect 119763 281931 119791 281959
rect 119577 281869 119605 281897
rect 119639 281869 119667 281897
rect 119701 281869 119729 281897
rect 119763 281869 119791 281897
rect 119577 281807 119605 281835
rect 119639 281807 119667 281835
rect 119701 281807 119729 281835
rect 119763 281807 119791 281835
rect 119577 281745 119605 281773
rect 119639 281745 119667 281773
rect 119701 281745 119729 281773
rect 119763 281745 119791 281773
rect 119577 272931 119605 272959
rect 119639 272931 119667 272959
rect 119701 272931 119729 272959
rect 119763 272931 119791 272959
rect 119577 272869 119605 272897
rect 119639 272869 119667 272897
rect 119701 272869 119729 272897
rect 119763 272869 119791 272897
rect 119577 272807 119605 272835
rect 119639 272807 119667 272835
rect 119701 272807 119729 272835
rect 119763 272807 119791 272835
rect 119577 272745 119605 272773
rect 119639 272745 119667 272773
rect 119701 272745 119729 272773
rect 119763 272745 119791 272773
rect 119577 263931 119605 263959
rect 119639 263931 119667 263959
rect 119701 263931 119729 263959
rect 119763 263931 119791 263959
rect 119577 263869 119605 263897
rect 119639 263869 119667 263897
rect 119701 263869 119729 263897
rect 119763 263869 119791 263897
rect 119577 263807 119605 263835
rect 119639 263807 119667 263835
rect 119701 263807 119729 263835
rect 119763 263807 119791 263835
rect 119577 263745 119605 263773
rect 119639 263745 119667 263773
rect 119701 263745 119729 263773
rect 119763 263745 119791 263773
rect 119577 254931 119605 254959
rect 119639 254931 119667 254959
rect 119701 254931 119729 254959
rect 119763 254931 119791 254959
rect 119577 254869 119605 254897
rect 119639 254869 119667 254897
rect 119701 254869 119729 254897
rect 119763 254869 119791 254897
rect 119577 254807 119605 254835
rect 119639 254807 119667 254835
rect 119701 254807 119729 254835
rect 119763 254807 119791 254835
rect 119577 254745 119605 254773
rect 119639 254745 119667 254773
rect 119701 254745 119729 254773
rect 119763 254745 119791 254773
rect 121437 299642 121465 299670
rect 121499 299642 121527 299670
rect 121561 299642 121589 299670
rect 121623 299642 121651 299670
rect 121437 299580 121465 299608
rect 121499 299580 121527 299608
rect 121561 299580 121589 299608
rect 121623 299580 121651 299608
rect 121437 299518 121465 299546
rect 121499 299518 121527 299546
rect 121561 299518 121589 299546
rect 121623 299518 121651 299546
rect 121437 299456 121465 299484
rect 121499 299456 121527 299484
rect 121561 299456 121589 299484
rect 121623 299456 121651 299484
rect 121437 293931 121465 293959
rect 121499 293931 121527 293959
rect 121561 293931 121589 293959
rect 121623 293931 121651 293959
rect 121437 293869 121465 293897
rect 121499 293869 121527 293897
rect 121561 293869 121589 293897
rect 121623 293869 121651 293897
rect 121437 293807 121465 293835
rect 121499 293807 121527 293835
rect 121561 293807 121589 293835
rect 121623 293807 121651 293835
rect 121437 293745 121465 293773
rect 121499 293745 121527 293773
rect 121561 293745 121589 293773
rect 121623 293745 121651 293773
rect 121437 284931 121465 284959
rect 121499 284931 121527 284959
rect 121561 284931 121589 284959
rect 121623 284931 121651 284959
rect 121437 284869 121465 284897
rect 121499 284869 121527 284897
rect 121561 284869 121589 284897
rect 121623 284869 121651 284897
rect 121437 284807 121465 284835
rect 121499 284807 121527 284835
rect 121561 284807 121589 284835
rect 121623 284807 121651 284835
rect 121437 284745 121465 284773
rect 121499 284745 121527 284773
rect 121561 284745 121589 284773
rect 121623 284745 121651 284773
rect 121437 275931 121465 275959
rect 121499 275931 121527 275959
rect 121561 275931 121589 275959
rect 121623 275931 121651 275959
rect 121437 275869 121465 275897
rect 121499 275869 121527 275897
rect 121561 275869 121589 275897
rect 121623 275869 121651 275897
rect 121437 275807 121465 275835
rect 121499 275807 121527 275835
rect 121561 275807 121589 275835
rect 121623 275807 121651 275835
rect 121437 275745 121465 275773
rect 121499 275745 121527 275773
rect 121561 275745 121589 275773
rect 121623 275745 121651 275773
rect 121437 266931 121465 266959
rect 121499 266931 121527 266959
rect 121561 266931 121589 266959
rect 121623 266931 121651 266959
rect 121437 266869 121465 266897
rect 121499 266869 121527 266897
rect 121561 266869 121589 266897
rect 121623 266869 121651 266897
rect 121437 266807 121465 266835
rect 121499 266807 121527 266835
rect 121561 266807 121589 266835
rect 121623 266807 121651 266835
rect 121437 266745 121465 266773
rect 121499 266745 121527 266773
rect 121561 266745 121589 266773
rect 121623 266745 121651 266773
rect 121437 257931 121465 257959
rect 121499 257931 121527 257959
rect 121561 257931 121589 257959
rect 121623 257931 121651 257959
rect 121437 257869 121465 257897
rect 121499 257869 121527 257897
rect 121561 257869 121589 257897
rect 121623 257869 121651 257897
rect 121437 257807 121465 257835
rect 121499 257807 121527 257835
rect 121561 257807 121589 257835
rect 121623 257807 121651 257835
rect 121437 257745 121465 257773
rect 121499 257745 121527 257773
rect 121561 257745 121589 257773
rect 121623 257745 121651 257773
rect 128577 299162 128605 299190
rect 128639 299162 128667 299190
rect 128701 299162 128729 299190
rect 128763 299162 128791 299190
rect 128577 299100 128605 299128
rect 128639 299100 128667 299128
rect 128701 299100 128729 299128
rect 128763 299100 128791 299128
rect 128577 299038 128605 299066
rect 128639 299038 128667 299066
rect 128701 299038 128729 299066
rect 128763 299038 128791 299066
rect 128577 298976 128605 299004
rect 128639 298976 128667 299004
rect 128701 298976 128729 299004
rect 128763 298976 128791 299004
rect 128577 290931 128605 290959
rect 128639 290931 128667 290959
rect 128701 290931 128729 290959
rect 128763 290931 128791 290959
rect 128577 290869 128605 290897
rect 128639 290869 128667 290897
rect 128701 290869 128729 290897
rect 128763 290869 128791 290897
rect 128577 290807 128605 290835
rect 128639 290807 128667 290835
rect 128701 290807 128729 290835
rect 128763 290807 128791 290835
rect 128577 290745 128605 290773
rect 128639 290745 128667 290773
rect 128701 290745 128729 290773
rect 128763 290745 128791 290773
rect 128577 281931 128605 281959
rect 128639 281931 128667 281959
rect 128701 281931 128729 281959
rect 128763 281931 128791 281959
rect 128577 281869 128605 281897
rect 128639 281869 128667 281897
rect 128701 281869 128729 281897
rect 128763 281869 128791 281897
rect 128577 281807 128605 281835
rect 128639 281807 128667 281835
rect 128701 281807 128729 281835
rect 128763 281807 128791 281835
rect 128577 281745 128605 281773
rect 128639 281745 128667 281773
rect 128701 281745 128729 281773
rect 128763 281745 128791 281773
rect 128577 272931 128605 272959
rect 128639 272931 128667 272959
rect 128701 272931 128729 272959
rect 128763 272931 128791 272959
rect 128577 272869 128605 272897
rect 128639 272869 128667 272897
rect 128701 272869 128729 272897
rect 128763 272869 128791 272897
rect 128577 272807 128605 272835
rect 128639 272807 128667 272835
rect 128701 272807 128729 272835
rect 128763 272807 128791 272835
rect 128577 272745 128605 272773
rect 128639 272745 128667 272773
rect 128701 272745 128729 272773
rect 128763 272745 128791 272773
rect 128577 263931 128605 263959
rect 128639 263931 128667 263959
rect 128701 263931 128729 263959
rect 128763 263931 128791 263959
rect 128577 263869 128605 263897
rect 128639 263869 128667 263897
rect 128701 263869 128729 263897
rect 128763 263869 128791 263897
rect 128577 263807 128605 263835
rect 128639 263807 128667 263835
rect 128701 263807 128729 263835
rect 128763 263807 128791 263835
rect 128577 263745 128605 263773
rect 128639 263745 128667 263773
rect 128701 263745 128729 263773
rect 128763 263745 128791 263773
rect 128577 254931 128605 254959
rect 128639 254931 128667 254959
rect 128701 254931 128729 254959
rect 128763 254931 128791 254959
rect 128577 254869 128605 254897
rect 128639 254869 128667 254897
rect 128701 254869 128729 254897
rect 128763 254869 128791 254897
rect 128577 254807 128605 254835
rect 128639 254807 128667 254835
rect 128701 254807 128729 254835
rect 128763 254807 128791 254835
rect 128577 254745 128605 254773
rect 128639 254745 128667 254773
rect 128701 254745 128729 254773
rect 128763 254745 128791 254773
rect 130437 299642 130465 299670
rect 130499 299642 130527 299670
rect 130561 299642 130589 299670
rect 130623 299642 130651 299670
rect 130437 299580 130465 299608
rect 130499 299580 130527 299608
rect 130561 299580 130589 299608
rect 130623 299580 130651 299608
rect 130437 299518 130465 299546
rect 130499 299518 130527 299546
rect 130561 299518 130589 299546
rect 130623 299518 130651 299546
rect 130437 299456 130465 299484
rect 130499 299456 130527 299484
rect 130561 299456 130589 299484
rect 130623 299456 130651 299484
rect 130437 293931 130465 293959
rect 130499 293931 130527 293959
rect 130561 293931 130589 293959
rect 130623 293931 130651 293959
rect 130437 293869 130465 293897
rect 130499 293869 130527 293897
rect 130561 293869 130589 293897
rect 130623 293869 130651 293897
rect 130437 293807 130465 293835
rect 130499 293807 130527 293835
rect 130561 293807 130589 293835
rect 130623 293807 130651 293835
rect 130437 293745 130465 293773
rect 130499 293745 130527 293773
rect 130561 293745 130589 293773
rect 130623 293745 130651 293773
rect 130437 284931 130465 284959
rect 130499 284931 130527 284959
rect 130561 284931 130589 284959
rect 130623 284931 130651 284959
rect 130437 284869 130465 284897
rect 130499 284869 130527 284897
rect 130561 284869 130589 284897
rect 130623 284869 130651 284897
rect 130437 284807 130465 284835
rect 130499 284807 130527 284835
rect 130561 284807 130589 284835
rect 130623 284807 130651 284835
rect 130437 284745 130465 284773
rect 130499 284745 130527 284773
rect 130561 284745 130589 284773
rect 130623 284745 130651 284773
rect 130437 275931 130465 275959
rect 130499 275931 130527 275959
rect 130561 275931 130589 275959
rect 130623 275931 130651 275959
rect 130437 275869 130465 275897
rect 130499 275869 130527 275897
rect 130561 275869 130589 275897
rect 130623 275869 130651 275897
rect 130437 275807 130465 275835
rect 130499 275807 130527 275835
rect 130561 275807 130589 275835
rect 130623 275807 130651 275835
rect 130437 275745 130465 275773
rect 130499 275745 130527 275773
rect 130561 275745 130589 275773
rect 130623 275745 130651 275773
rect 130437 266931 130465 266959
rect 130499 266931 130527 266959
rect 130561 266931 130589 266959
rect 130623 266931 130651 266959
rect 130437 266869 130465 266897
rect 130499 266869 130527 266897
rect 130561 266869 130589 266897
rect 130623 266869 130651 266897
rect 130437 266807 130465 266835
rect 130499 266807 130527 266835
rect 130561 266807 130589 266835
rect 130623 266807 130651 266835
rect 130437 266745 130465 266773
rect 130499 266745 130527 266773
rect 130561 266745 130589 266773
rect 130623 266745 130651 266773
rect 130437 257931 130465 257959
rect 130499 257931 130527 257959
rect 130561 257931 130589 257959
rect 130623 257931 130651 257959
rect 130437 257869 130465 257897
rect 130499 257869 130527 257897
rect 130561 257869 130589 257897
rect 130623 257869 130651 257897
rect 130437 257807 130465 257835
rect 130499 257807 130527 257835
rect 130561 257807 130589 257835
rect 130623 257807 130651 257835
rect 130437 257745 130465 257773
rect 130499 257745 130527 257773
rect 130561 257745 130589 257773
rect 130623 257745 130651 257773
rect 137577 299162 137605 299190
rect 137639 299162 137667 299190
rect 137701 299162 137729 299190
rect 137763 299162 137791 299190
rect 137577 299100 137605 299128
rect 137639 299100 137667 299128
rect 137701 299100 137729 299128
rect 137763 299100 137791 299128
rect 137577 299038 137605 299066
rect 137639 299038 137667 299066
rect 137701 299038 137729 299066
rect 137763 299038 137791 299066
rect 137577 298976 137605 299004
rect 137639 298976 137667 299004
rect 137701 298976 137729 299004
rect 137763 298976 137791 299004
rect 137577 290931 137605 290959
rect 137639 290931 137667 290959
rect 137701 290931 137729 290959
rect 137763 290931 137791 290959
rect 137577 290869 137605 290897
rect 137639 290869 137667 290897
rect 137701 290869 137729 290897
rect 137763 290869 137791 290897
rect 137577 290807 137605 290835
rect 137639 290807 137667 290835
rect 137701 290807 137729 290835
rect 137763 290807 137791 290835
rect 137577 290745 137605 290773
rect 137639 290745 137667 290773
rect 137701 290745 137729 290773
rect 137763 290745 137791 290773
rect 137577 281931 137605 281959
rect 137639 281931 137667 281959
rect 137701 281931 137729 281959
rect 137763 281931 137791 281959
rect 137577 281869 137605 281897
rect 137639 281869 137667 281897
rect 137701 281869 137729 281897
rect 137763 281869 137791 281897
rect 137577 281807 137605 281835
rect 137639 281807 137667 281835
rect 137701 281807 137729 281835
rect 137763 281807 137791 281835
rect 137577 281745 137605 281773
rect 137639 281745 137667 281773
rect 137701 281745 137729 281773
rect 137763 281745 137791 281773
rect 137577 272931 137605 272959
rect 137639 272931 137667 272959
rect 137701 272931 137729 272959
rect 137763 272931 137791 272959
rect 137577 272869 137605 272897
rect 137639 272869 137667 272897
rect 137701 272869 137729 272897
rect 137763 272869 137791 272897
rect 137577 272807 137605 272835
rect 137639 272807 137667 272835
rect 137701 272807 137729 272835
rect 137763 272807 137791 272835
rect 137577 272745 137605 272773
rect 137639 272745 137667 272773
rect 137701 272745 137729 272773
rect 137763 272745 137791 272773
rect 137577 263931 137605 263959
rect 137639 263931 137667 263959
rect 137701 263931 137729 263959
rect 137763 263931 137791 263959
rect 137577 263869 137605 263897
rect 137639 263869 137667 263897
rect 137701 263869 137729 263897
rect 137763 263869 137791 263897
rect 137577 263807 137605 263835
rect 137639 263807 137667 263835
rect 137701 263807 137729 263835
rect 137763 263807 137791 263835
rect 137577 263745 137605 263773
rect 137639 263745 137667 263773
rect 137701 263745 137729 263773
rect 137763 263745 137791 263773
rect 137577 254931 137605 254959
rect 137639 254931 137667 254959
rect 137701 254931 137729 254959
rect 137763 254931 137791 254959
rect 137577 254869 137605 254897
rect 137639 254869 137667 254897
rect 137701 254869 137729 254897
rect 137763 254869 137791 254897
rect 137577 254807 137605 254835
rect 137639 254807 137667 254835
rect 137701 254807 137729 254835
rect 137763 254807 137791 254835
rect 137577 254745 137605 254773
rect 137639 254745 137667 254773
rect 137701 254745 137729 254773
rect 137763 254745 137791 254773
rect 139437 299642 139465 299670
rect 139499 299642 139527 299670
rect 139561 299642 139589 299670
rect 139623 299642 139651 299670
rect 139437 299580 139465 299608
rect 139499 299580 139527 299608
rect 139561 299580 139589 299608
rect 139623 299580 139651 299608
rect 139437 299518 139465 299546
rect 139499 299518 139527 299546
rect 139561 299518 139589 299546
rect 139623 299518 139651 299546
rect 139437 299456 139465 299484
rect 139499 299456 139527 299484
rect 139561 299456 139589 299484
rect 139623 299456 139651 299484
rect 139437 293931 139465 293959
rect 139499 293931 139527 293959
rect 139561 293931 139589 293959
rect 139623 293931 139651 293959
rect 139437 293869 139465 293897
rect 139499 293869 139527 293897
rect 139561 293869 139589 293897
rect 139623 293869 139651 293897
rect 139437 293807 139465 293835
rect 139499 293807 139527 293835
rect 139561 293807 139589 293835
rect 139623 293807 139651 293835
rect 139437 293745 139465 293773
rect 139499 293745 139527 293773
rect 139561 293745 139589 293773
rect 139623 293745 139651 293773
rect 139437 284931 139465 284959
rect 139499 284931 139527 284959
rect 139561 284931 139589 284959
rect 139623 284931 139651 284959
rect 139437 284869 139465 284897
rect 139499 284869 139527 284897
rect 139561 284869 139589 284897
rect 139623 284869 139651 284897
rect 139437 284807 139465 284835
rect 139499 284807 139527 284835
rect 139561 284807 139589 284835
rect 139623 284807 139651 284835
rect 139437 284745 139465 284773
rect 139499 284745 139527 284773
rect 139561 284745 139589 284773
rect 139623 284745 139651 284773
rect 139437 275931 139465 275959
rect 139499 275931 139527 275959
rect 139561 275931 139589 275959
rect 139623 275931 139651 275959
rect 139437 275869 139465 275897
rect 139499 275869 139527 275897
rect 139561 275869 139589 275897
rect 139623 275869 139651 275897
rect 139437 275807 139465 275835
rect 139499 275807 139527 275835
rect 139561 275807 139589 275835
rect 139623 275807 139651 275835
rect 139437 275745 139465 275773
rect 139499 275745 139527 275773
rect 139561 275745 139589 275773
rect 139623 275745 139651 275773
rect 139437 266931 139465 266959
rect 139499 266931 139527 266959
rect 139561 266931 139589 266959
rect 139623 266931 139651 266959
rect 139437 266869 139465 266897
rect 139499 266869 139527 266897
rect 139561 266869 139589 266897
rect 139623 266869 139651 266897
rect 139437 266807 139465 266835
rect 139499 266807 139527 266835
rect 139561 266807 139589 266835
rect 139623 266807 139651 266835
rect 139437 266745 139465 266773
rect 139499 266745 139527 266773
rect 139561 266745 139589 266773
rect 139623 266745 139651 266773
rect 139437 257931 139465 257959
rect 139499 257931 139527 257959
rect 139561 257931 139589 257959
rect 139623 257931 139651 257959
rect 139437 257869 139465 257897
rect 139499 257869 139527 257897
rect 139561 257869 139589 257897
rect 139623 257869 139651 257897
rect 139437 257807 139465 257835
rect 139499 257807 139527 257835
rect 139561 257807 139589 257835
rect 139623 257807 139651 257835
rect 139437 257745 139465 257773
rect 139499 257745 139527 257773
rect 139561 257745 139589 257773
rect 139623 257745 139651 257773
rect 146577 299162 146605 299190
rect 146639 299162 146667 299190
rect 146701 299162 146729 299190
rect 146763 299162 146791 299190
rect 146577 299100 146605 299128
rect 146639 299100 146667 299128
rect 146701 299100 146729 299128
rect 146763 299100 146791 299128
rect 146577 299038 146605 299066
rect 146639 299038 146667 299066
rect 146701 299038 146729 299066
rect 146763 299038 146791 299066
rect 146577 298976 146605 299004
rect 146639 298976 146667 299004
rect 146701 298976 146729 299004
rect 146763 298976 146791 299004
rect 146577 290931 146605 290959
rect 146639 290931 146667 290959
rect 146701 290931 146729 290959
rect 146763 290931 146791 290959
rect 146577 290869 146605 290897
rect 146639 290869 146667 290897
rect 146701 290869 146729 290897
rect 146763 290869 146791 290897
rect 146577 290807 146605 290835
rect 146639 290807 146667 290835
rect 146701 290807 146729 290835
rect 146763 290807 146791 290835
rect 146577 290745 146605 290773
rect 146639 290745 146667 290773
rect 146701 290745 146729 290773
rect 146763 290745 146791 290773
rect 146577 281931 146605 281959
rect 146639 281931 146667 281959
rect 146701 281931 146729 281959
rect 146763 281931 146791 281959
rect 146577 281869 146605 281897
rect 146639 281869 146667 281897
rect 146701 281869 146729 281897
rect 146763 281869 146791 281897
rect 146577 281807 146605 281835
rect 146639 281807 146667 281835
rect 146701 281807 146729 281835
rect 146763 281807 146791 281835
rect 146577 281745 146605 281773
rect 146639 281745 146667 281773
rect 146701 281745 146729 281773
rect 146763 281745 146791 281773
rect 146577 272931 146605 272959
rect 146639 272931 146667 272959
rect 146701 272931 146729 272959
rect 146763 272931 146791 272959
rect 146577 272869 146605 272897
rect 146639 272869 146667 272897
rect 146701 272869 146729 272897
rect 146763 272869 146791 272897
rect 146577 272807 146605 272835
rect 146639 272807 146667 272835
rect 146701 272807 146729 272835
rect 146763 272807 146791 272835
rect 146577 272745 146605 272773
rect 146639 272745 146667 272773
rect 146701 272745 146729 272773
rect 146763 272745 146791 272773
rect 146577 263931 146605 263959
rect 146639 263931 146667 263959
rect 146701 263931 146729 263959
rect 146763 263931 146791 263959
rect 146577 263869 146605 263897
rect 146639 263869 146667 263897
rect 146701 263869 146729 263897
rect 146763 263869 146791 263897
rect 146577 263807 146605 263835
rect 146639 263807 146667 263835
rect 146701 263807 146729 263835
rect 146763 263807 146791 263835
rect 146577 263745 146605 263773
rect 146639 263745 146667 263773
rect 146701 263745 146729 263773
rect 146763 263745 146791 263773
rect 146577 254931 146605 254959
rect 146639 254931 146667 254959
rect 146701 254931 146729 254959
rect 146763 254931 146791 254959
rect 146577 254869 146605 254897
rect 146639 254869 146667 254897
rect 146701 254869 146729 254897
rect 146763 254869 146791 254897
rect 146577 254807 146605 254835
rect 146639 254807 146667 254835
rect 146701 254807 146729 254835
rect 146763 254807 146791 254835
rect 146577 254745 146605 254773
rect 146639 254745 146667 254773
rect 146701 254745 146729 254773
rect 146763 254745 146791 254773
rect 148437 299642 148465 299670
rect 148499 299642 148527 299670
rect 148561 299642 148589 299670
rect 148623 299642 148651 299670
rect 148437 299580 148465 299608
rect 148499 299580 148527 299608
rect 148561 299580 148589 299608
rect 148623 299580 148651 299608
rect 148437 299518 148465 299546
rect 148499 299518 148527 299546
rect 148561 299518 148589 299546
rect 148623 299518 148651 299546
rect 148437 299456 148465 299484
rect 148499 299456 148527 299484
rect 148561 299456 148589 299484
rect 148623 299456 148651 299484
rect 148437 293931 148465 293959
rect 148499 293931 148527 293959
rect 148561 293931 148589 293959
rect 148623 293931 148651 293959
rect 148437 293869 148465 293897
rect 148499 293869 148527 293897
rect 148561 293869 148589 293897
rect 148623 293869 148651 293897
rect 148437 293807 148465 293835
rect 148499 293807 148527 293835
rect 148561 293807 148589 293835
rect 148623 293807 148651 293835
rect 148437 293745 148465 293773
rect 148499 293745 148527 293773
rect 148561 293745 148589 293773
rect 148623 293745 148651 293773
rect 148437 284931 148465 284959
rect 148499 284931 148527 284959
rect 148561 284931 148589 284959
rect 148623 284931 148651 284959
rect 148437 284869 148465 284897
rect 148499 284869 148527 284897
rect 148561 284869 148589 284897
rect 148623 284869 148651 284897
rect 148437 284807 148465 284835
rect 148499 284807 148527 284835
rect 148561 284807 148589 284835
rect 148623 284807 148651 284835
rect 148437 284745 148465 284773
rect 148499 284745 148527 284773
rect 148561 284745 148589 284773
rect 148623 284745 148651 284773
rect 148437 275931 148465 275959
rect 148499 275931 148527 275959
rect 148561 275931 148589 275959
rect 148623 275931 148651 275959
rect 148437 275869 148465 275897
rect 148499 275869 148527 275897
rect 148561 275869 148589 275897
rect 148623 275869 148651 275897
rect 148437 275807 148465 275835
rect 148499 275807 148527 275835
rect 148561 275807 148589 275835
rect 148623 275807 148651 275835
rect 148437 275745 148465 275773
rect 148499 275745 148527 275773
rect 148561 275745 148589 275773
rect 148623 275745 148651 275773
rect 148437 266931 148465 266959
rect 148499 266931 148527 266959
rect 148561 266931 148589 266959
rect 148623 266931 148651 266959
rect 148437 266869 148465 266897
rect 148499 266869 148527 266897
rect 148561 266869 148589 266897
rect 148623 266869 148651 266897
rect 148437 266807 148465 266835
rect 148499 266807 148527 266835
rect 148561 266807 148589 266835
rect 148623 266807 148651 266835
rect 148437 266745 148465 266773
rect 148499 266745 148527 266773
rect 148561 266745 148589 266773
rect 148623 266745 148651 266773
rect 148437 257931 148465 257959
rect 148499 257931 148527 257959
rect 148561 257931 148589 257959
rect 148623 257931 148651 257959
rect 148437 257869 148465 257897
rect 148499 257869 148527 257897
rect 148561 257869 148589 257897
rect 148623 257869 148651 257897
rect 148437 257807 148465 257835
rect 148499 257807 148527 257835
rect 148561 257807 148589 257835
rect 148623 257807 148651 257835
rect 148437 257745 148465 257773
rect 148499 257745 148527 257773
rect 148561 257745 148589 257773
rect 148623 257745 148651 257773
rect 155577 299162 155605 299190
rect 155639 299162 155667 299190
rect 155701 299162 155729 299190
rect 155763 299162 155791 299190
rect 155577 299100 155605 299128
rect 155639 299100 155667 299128
rect 155701 299100 155729 299128
rect 155763 299100 155791 299128
rect 155577 299038 155605 299066
rect 155639 299038 155667 299066
rect 155701 299038 155729 299066
rect 155763 299038 155791 299066
rect 155577 298976 155605 299004
rect 155639 298976 155667 299004
rect 155701 298976 155729 299004
rect 155763 298976 155791 299004
rect 155577 290931 155605 290959
rect 155639 290931 155667 290959
rect 155701 290931 155729 290959
rect 155763 290931 155791 290959
rect 155577 290869 155605 290897
rect 155639 290869 155667 290897
rect 155701 290869 155729 290897
rect 155763 290869 155791 290897
rect 155577 290807 155605 290835
rect 155639 290807 155667 290835
rect 155701 290807 155729 290835
rect 155763 290807 155791 290835
rect 155577 290745 155605 290773
rect 155639 290745 155667 290773
rect 155701 290745 155729 290773
rect 155763 290745 155791 290773
rect 155577 281931 155605 281959
rect 155639 281931 155667 281959
rect 155701 281931 155729 281959
rect 155763 281931 155791 281959
rect 155577 281869 155605 281897
rect 155639 281869 155667 281897
rect 155701 281869 155729 281897
rect 155763 281869 155791 281897
rect 155577 281807 155605 281835
rect 155639 281807 155667 281835
rect 155701 281807 155729 281835
rect 155763 281807 155791 281835
rect 155577 281745 155605 281773
rect 155639 281745 155667 281773
rect 155701 281745 155729 281773
rect 155763 281745 155791 281773
rect 155577 272931 155605 272959
rect 155639 272931 155667 272959
rect 155701 272931 155729 272959
rect 155763 272931 155791 272959
rect 155577 272869 155605 272897
rect 155639 272869 155667 272897
rect 155701 272869 155729 272897
rect 155763 272869 155791 272897
rect 155577 272807 155605 272835
rect 155639 272807 155667 272835
rect 155701 272807 155729 272835
rect 155763 272807 155791 272835
rect 155577 272745 155605 272773
rect 155639 272745 155667 272773
rect 155701 272745 155729 272773
rect 155763 272745 155791 272773
rect 155577 263931 155605 263959
rect 155639 263931 155667 263959
rect 155701 263931 155729 263959
rect 155763 263931 155791 263959
rect 155577 263869 155605 263897
rect 155639 263869 155667 263897
rect 155701 263869 155729 263897
rect 155763 263869 155791 263897
rect 155577 263807 155605 263835
rect 155639 263807 155667 263835
rect 155701 263807 155729 263835
rect 155763 263807 155791 263835
rect 155577 263745 155605 263773
rect 155639 263745 155667 263773
rect 155701 263745 155729 263773
rect 155763 263745 155791 263773
rect 155577 254931 155605 254959
rect 155639 254931 155667 254959
rect 155701 254931 155729 254959
rect 155763 254931 155791 254959
rect 155577 254869 155605 254897
rect 155639 254869 155667 254897
rect 155701 254869 155729 254897
rect 155763 254869 155791 254897
rect 155577 254807 155605 254835
rect 155639 254807 155667 254835
rect 155701 254807 155729 254835
rect 155763 254807 155791 254835
rect 155577 254745 155605 254773
rect 155639 254745 155667 254773
rect 155701 254745 155729 254773
rect 155763 254745 155791 254773
rect 157437 299642 157465 299670
rect 157499 299642 157527 299670
rect 157561 299642 157589 299670
rect 157623 299642 157651 299670
rect 157437 299580 157465 299608
rect 157499 299580 157527 299608
rect 157561 299580 157589 299608
rect 157623 299580 157651 299608
rect 157437 299518 157465 299546
rect 157499 299518 157527 299546
rect 157561 299518 157589 299546
rect 157623 299518 157651 299546
rect 157437 299456 157465 299484
rect 157499 299456 157527 299484
rect 157561 299456 157589 299484
rect 157623 299456 157651 299484
rect 157437 293931 157465 293959
rect 157499 293931 157527 293959
rect 157561 293931 157589 293959
rect 157623 293931 157651 293959
rect 157437 293869 157465 293897
rect 157499 293869 157527 293897
rect 157561 293869 157589 293897
rect 157623 293869 157651 293897
rect 157437 293807 157465 293835
rect 157499 293807 157527 293835
rect 157561 293807 157589 293835
rect 157623 293807 157651 293835
rect 157437 293745 157465 293773
rect 157499 293745 157527 293773
rect 157561 293745 157589 293773
rect 157623 293745 157651 293773
rect 157437 284931 157465 284959
rect 157499 284931 157527 284959
rect 157561 284931 157589 284959
rect 157623 284931 157651 284959
rect 157437 284869 157465 284897
rect 157499 284869 157527 284897
rect 157561 284869 157589 284897
rect 157623 284869 157651 284897
rect 157437 284807 157465 284835
rect 157499 284807 157527 284835
rect 157561 284807 157589 284835
rect 157623 284807 157651 284835
rect 157437 284745 157465 284773
rect 157499 284745 157527 284773
rect 157561 284745 157589 284773
rect 157623 284745 157651 284773
rect 157437 275931 157465 275959
rect 157499 275931 157527 275959
rect 157561 275931 157589 275959
rect 157623 275931 157651 275959
rect 157437 275869 157465 275897
rect 157499 275869 157527 275897
rect 157561 275869 157589 275897
rect 157623 275869 157651 275897
rect 157437 275807 157465 275835
rect 157499 275807 157527 275835
rect 157561 275807 157589 275835
rect 157623 275807 157651 275835
rect 157437 275745 157465 275773
rect 157499 275745 157527 275773
rect 157561 275745 157589 275773
rect 157623 275745 157651 275773
rect 157437 266931 157465 266959
rect 157499 266931 157527 266959
rect 157561 266931 157589 266959
rect 157623 266931 157651 266959
rect 157437 266869 157465 266897
rect 157499 266869 157527 266897
rect 157561 266869 157589 266897
rect 157623 266869 157651 266897
rect 157437 266807 157465 266835
rect 157499 266807 157527 266835
rect 157561 266807 157589 266835
rect 157623 266807 157651 266835
rect 157437 266745 157465 266773
rect 157499 266745 157527 266773
rect 157561 266745 157589 266773
rect 157623 266745 157651 266773
rect 157437 257931 157465 257959
rect 157499 257931 157527 257959
rect 157561 257931 157589 257959
rect 157623 257931 157651 257959
rect 157437 257869 157465 257897
rect 157499 257869 157527 257897
rect 157561 257869 157589 257897
rect 157623 257869 157651 257897
rect 157437 257807 157465 257835
rect 157499 257807 157527 257835
rect 157561 257807 157589 257835
rect 157623 257807 157651 257835
rect 157437 257745 157465 257773
rect 157499 257745 157527 257773
rect 157561 257745 157589 257773
rect 157623 257745 157651 257773
rect 164577 299162 164605 299190
rect 164639 299162 164667 299190
rect 164701 299162 164729 299190
rect 164763 299162 164791 299190
rect 164577 299100 164605 299128
rect 164639 299100 164667 299128
rect 164701 299100 164729 299128
rect 164763 299100 164791 299128
rect 164577 299038 164605 299066
rect 164639 299038 164667 299066
rect 164701 299038 164729 299066
rect 164763 299038 164791 299066
rect 164577 298976 164605 299004
rect 164639 298976 164667 299004
rect 164701 298976 164729 299004
rect 164763 298976 164791 299004
rect 164577 290931 164605 290959
rect 164639 290931 164667 290959
rect 164701 290931 164729 290959
rect 164763 290931 164791 290959
rect 164577 290869 164605 290897
rect 164639 290869 164667 290897
rect 164701 290869 164729 290897
rect 164763 290869 164791 290897
rect 164577 290807 164605 290835
rect 164639 290807 164667 290835
rect 164701 290807 164729 290835
rect 164763 290807 164791 290835
rect 164577 290745 164605 290773
rect 164639 290745 164667 290773
rect 164701 290745 164729 290773
rect 164763 290745 164791 290773
rect 164577 281931 164605 281959
rect 164639 281931 164667 281959
rect 164701 281931 164729 281959
rect 164763 281931 164791 281959
rect 164577 281869 164605 281897
rect 164639 281869 164667 281897
rect 164701 281869 164729 281897
rect 164763 281869 164791 281897
rect 164577 281807 164605 281835
rect 164639 281807 164667 281835
rect 164701 281807 164729 281835
rect 164763 281807 164791 281835
rect 164577 281745 164605 281773
rect 164639 281745 164667 281773
rect 164701 281745 164729 281773
rect 164763 281745 164791 281773
rect 164577 272931 164605 272959
rect 164639 272931 164667 272959
rect 164701 272931 164729 272959
rect 164763 272931 164791 272959
rect 164577 272869 164605 272897
rect 164639 272869 164667 272897
rect 164701 272869 164729 272897
rect 164763 272869 164791 272897
rect 164577 272807 164605 272835
rect 164639 272807 164667 272835
rect 164701 272807 164729 272835
rect 164763 272807 164791 272835
rect 164577 272745 164605 272773
rect 164639 272745 164667 272773
rect 164701 272745 164729 272773
rect 164763 272745 164791 272773
rect 164577 263931 164605 263959
rect 164639 263931 164667 263959
rect 164701 263931 164729 263959
rect 164763 263931 164791 263959
rect 164577 263869 164605 263897
rect 164639 263869 164667 263897
rect 164701 263869 164729 263897
rect 164763 263869 164791 263897
rect 164577 263807 164605 263835
rect 164639 263807 164667 263835
rect 164701 263807 164729 263835
rect 164763 263807 164791 263835
rect 164577 263745 164605 263773
rect 164639 263745 164667 263773
rect 164701 263745 164729 263773
rect 164763 263745 164791 263773
rect 164577 254931 164605 254959
rect 164639 254931 164667 254959
rect 164701 254931 164729 254959
rect 164763 254931 164791 254959
rect 164577 254869 164605 254897
rect 164639 254869 164667 254897
rect 164701 254869 164729 254897
rect 164763 254869 164791 254897
rect 164577 254807 164605 254835
rect 164639 254807 164667 254835
rect 164701 254807 164729 254835
rect 164763 254807 164791 254835
rect 164577 254745 164605 254773
rect 164639 254745 164667 254773
rect 164701 254745 164729 254773
rect 164763 254745 164791 254773
rect 166437 299642 166465 299670
rect 166499 299642 166527 299670
rect 166561 299642 166589 299670
rect 166623 299642 166651 299670
rect 166437 299580 166465 299608
rect 166499 299580 166527 299608
rect 166561 299580 166589 299608
rect 166623 299580 166651 299608
rect 166437 299518 166465 299546
rect 166499 299518 166527 299546
rect 166561 299518 166589 299546
rect 166623 299518 166651 299546
rect 166437 299456 166465 299484
rect 166499 299456 166527 299484
rect 166561 299456 166589 299484
rect 166623 299456 166651 299484
rect 166437 293931 166465 293959
rect 166499 293931 166527 293959
rect 166561 293931 166589 293959
rect 166623 293931 166651 293959
rect 166437 293869 166465 293897
rect 166499 293869 166527 293897
rect 166561 293869 166589 293897
rect 166623 293869 166651 293897
rect 166437 293807 166465 293835
rect 166499 293807 166527 293835
rect 166561 293807 166589 293835
rect 166623 293807 166651 293835
rect 166437 293745 166465 293773
rect 166499 293745 166527 293773
rect 166561 293745 166589 293773
rect 166623 293745 166651 293773
rect 166437 284931 166465 284959
rect 166499 284931 166527 284959
rect 166561 284931 166589 284959
rect 166623 284931 166651 284959
rect 166437 284869 166465 284897
rect 166499 284869 166527 284897
rect 166561 284869 166589 284897
rect 166623 284869 166651 284897
rect 166437 284807 166465 284835
rect 166499 284807 166527 284835
rect 166561 284807 166589 284835
rect 166623 284807 166651 284835
rect 166437 284745 166465 284773
rect 166499 284745 166527 284773
rect 166561 284745 166589 284773
rect 166623 284745 166651 284773
rect 166437 275931 166465 275959
rect 166499 275931 166527 275959
rect 166561 275931 166589 275959
rect 166623 275931 166651 275959
rect 166437 275869 166465 275897
rect 166499 275869 166527 275897
rect 166561 275869 166589 275897
rect 166623 275869 166651 275897
rect 166437 275807 166465 275835
rect 166499 275807 166527 275835
rect 166561 275807 166589 275835
rect 166623 275807 166651 275835
rect 166437 275745 166465 275773
rect 166499 275745 166527 275773
rect 166561 275745 166589 275773
rect 166623 275745 166651 275773
rect 166437 266931 166465 266959
rect 166499 266931 166527 266959
rect 166561 266931 166589 266959
rect 166623 266931 166651 266959
rect 166437 266869 166465 266897
rect 166499 266869 166527 266897
rect 166561 266869 166589 266897
rect 166623 266869 166651 266897
rect 166437 266807 166465 266835
rect 166499 266807 166527 266835
rect 166561 266807 166589 266835
rect 166623 266807 166651 266835
rect 166437 266745 166465 266773
rect 166499 266745 166527 266773
rect 166561 266745 166589 266773
rect 166623 266745 166651 266773
rect 166437 257931 166465 257959
rect 166499 257931 166527 257959
rect 166561 257931 166589 257959
rect 166623 257931 166651 257959
rect 166437 257869 166465 257897
rect 166499 257869 166527 257897
rect 166561 257869 166589 257897
rect 166623 257869 166651 257897
rect 166437 257807 166465 257835
rect 166499 257807 166527 257835
rect 166561 257807 166589 257835
rect 166623 257807 166651 257835
rect 166437 257745 166465 257773
rect 166499 257745 166527 257773
rect 166561 257745 166589 257773
rect 166623 257745 166651 257773
rect 173577 299162 173605 299190
rect 173639 299162 173667 299190
rect 173701 299162 173729 299190
rect 173763 299162 173791 299190
rect 173577 299100 173605 299128
rect 173639 299100 173667 299128
rect 173701 299100 173729 299128
rect 173763 299100 173791 299128
rect 173577 299038 173605 299066
rect 173639 299038 173667 299066
rect 173701 299038 173729 299066
rect 173763 299038 173791 299066
rect 173577 298976 173605 299004
rect 173639 298976 173667 299004
rect 173701 298976 173729 299004
rect 173763 298976 173791 299004
rect 173577 290931 173605 290959
rect 173639 290931 173667 290959
rect 173701 290931 173729 290959
rect 173763 290931 173791 290959
rect 173577 290869 173605 290897
rect 173639 290869 173667 290897
rect 173701 290869 173729 290897
rect 173763 290869 173791 290897
rect 173577 290807 173605 290835
rect 173639 290807 173667 290835
rect 173701 290807 173729 290835
rect 173763 290807 173791 290835
rect 173577 290745 173605 290773
rect 173639 290745 173667 290773
rect 173701 290745 173729 290773
rect 173763 290745 173791 290773
rect 173577 281931 173605 281959
rect 173639 281931 173667 281959
rect 173701 281931 173729 281959
rect 173763 281931 173791 281959
rect 173577 281869 173605 281897
rect 173639 281869 173667 281897
rect 173701 281869 173729 281897
rect 173763 281869 173791 281897
rect 173577 281807 173605 281835
rect 173639 281807 173667 281835
rect 173701 281807 173729 281835
rect 173763 281807 173791 281835
rect 173577 281745 173605 281773
rect 173639 281745 173667 281773
rect 173701 281745 173729 281773
rect 173763 281745 173791 281773
rect 173577 272931 173605 272959
rect 173639 272931 173667 272959
rect 173701 272931 173729 272959
rect 173763 272931 173791 272959
rect 173577 272869 173605 272897
rect 173639 272869 173667 272897
rect 173701 272869 173729 272897
rect 173763 272869 173791 272897
rect 173577 272807 173605 272835
rect 173639 272807 173667 272835
rect 173701 272807 173729 272835
rect 173763 272807 173791 272835
rect 173577 272745 173605 272773
rect 173639 272745 173667 272773
rect 173701 272745 173729 272773
rect 173763 272745 173791 272773
rect 173577 263931 173605 263959
rect 173639 263931 173667 263959
rect 173701 263931 173729 263959
rect 173763 263931 173791 263959
rect 173577 263869 173605 263897
rect 173639 263869 173667 263897
rect 173701 263869 173729 263897
rect 173763 263869 173791 263897
rect 173577 263807 173605 263835
rect 173639 263807 173667 263835
rect 173701 263807 173729 263835
rect 173763 263807 173791 263835
rect 173577 263745 173605 263773
rect 173639 263745 173667 263773
rect 173701 263745 173729 263773
rect 173763 263745 173791 263773
rect 173577 254931 173605 254959
rect 173639 254931 173667 254959
rect 173701 254931 173729 254959
rect 173763 254931 173791 254959
rect 173577 254869 173605 254897
rect 173639 254869 173667 254897
rect 173701 254869 173729 254897
rect 173763 254869 173791 254897
rect 173577 254807 173605 254835
rect 173639 254807 173667 254835
rect 173701 254807 173729 254835
rect 173763 254807 173791 254835
rect 173577 254745 173605 254773
rect 173639 254745 173667 254773
rect 173701 254745 173729 254773
rect 173763 254745 173791 254773
rect 175437 299642 175465 299670
rect 175499 299642 175527 299670
rect 175561 299642 175589 299670
rect 175623 299642 175651 299670
rect 175437 299580 175465 299608
rect 175499 299580 175527 299608
rect 175561 299580 175589 299608
rect 175623 299580 175651 299608
rect 175437 299518 175465 299546
rect 175499 299518 175527 299546
rect 175561 299518 175589 299546
rect 175623 299518 175651 299546
rect 175437 299456 175465 299484
rect 175499 299456 175527 299484
rect 175561 299456 175589 299484
rect 175623 299456 175651 299484
rect 175437 293931 175465 293959
rect 175499 293931 175527 293959
rect 175561 293931 175589 293959
rect 175623 293931 175651 293959
rect 175437 293869 175465 293897
rect 175499 293869 175527 293897
rect 175561 293869 175589 293897
rect 175623 293869 175651 293897
rect 175437 293807 175465 293835
rect 175499 293807 175527 293835
rect 175561 293807 175589 293835
rect 175623 293807 175651 293835
rect 175437 293745 175465 293773
rect 175499 293745 175527 293773
rect 175561 293745 175589 293773
rect 175623 293745 175651 293773
rect 175437 284931 175465 284959
rect 175499 284931 175527 284959
rect 175561 284931 175589 284959
rect 175623 284931 175651 284959
rect 175437 284869 175465 284897
rect 175499 284869 175527 284897
rect 175561 284869 175589 284897
rect 175623 284869 175651 284897
rect 175437 284807 175465 284835
rect 175499 284807 175527 284835
rect 175561 284807 175589 284835
rect 175623 284807 175651 284835
rect 175437 284745 175465 284773
rect 175499 284745 175527 284773
rect 175561 284745 175589 284773
rect 175623 284745 175651 284773
rect 175437 275931 175465 275959
rect 175499 275931 175527 275959
rect 175561 275931 175589 275959
rect 175623 275931 175651 275959
rect 175437 275869 175465 275897
rect 175499 275869 175527 275897
rect 175561 275869 175589 275897
rect 175623 275869 175651 275897
rect 175437 275807 175465 275835
rect 175499 275807 175527 275835
rect 175561 275807 175589 275835
rect 175623 275807 175651 275835
rect 175437 275745 175465 275773
rect 175499 275745 175527 275773
rect 175561 275745 175589 275773
rect 175623 275745 175651 275773
rect 175437 266931 175465 266959
rect 175499 266931 175527 266959
rect 175561 266931 175589 266959
rect 175623 266931 175651 266959
rect 175437 266869 175465 266897
rect 175499 266869 175527 266897
rect 175561 266869 175589 266897
rect 175623 266869 175651 266897
rect 175437 266807 175465 266835
rect 175499 266807 175527 266835
rect 175561 266807 175589 266835
rect 175623 266807 175651 266835
rect 175437 266745 175465 266773
rect 175499 266745 175527 266773
rect 175561 266745 175589 266773
rect 175623 266745 175651 266773
rect 175437 257931 175465 257959
rect 175499 257931 175527 257959
rect 175561 257931 175589 257959
rect 175623 257931 175651 257959
rect 175437 257869 175465 257897
rect 175499 257869 175527 257897
rect 175561 257869 175589 257897
rect 175623 257869 175651 257897
rect 175437 257807 175465 257835
rect 175499 257807 175527 257835
rect 175561 257807 175589 257835
rect 175623 257807 175651 257835
rect 175437 257745 175465 257773
rect 175499 257745 175527 257773
rect 175561 257745 175589 257773
rect 175623 257745 175651 257773
rect 182577 299162 182605 299190
rect 182639 299162 182667 299190
rect 182701 299162 182729 299190
rect 182763 299162 182791 299190
rect 182577 299100 182605 299128
rect 182639 299100 182667 299128
rect 182701 299100 182729 299128
rect 182763 299100 182791 299128
rect 182577 299038 182605 299066
rect 182639 299038 182667 299066
rect 182701 299038 182729 299066
rect 182763 299038 182791 299066
rect 182577 298976 182605 299004
rect 182639 298976 182667 299004
rect 182701 298976 182729 299004
rect 182763 298976 182791 299004
rect 182577 290931 182605 290959
rect 182639 290931 182667 290959
rect 182701 290931 182729 290959
rect 182763 290931 182791 290959
rect 182577 290869 182605 290897
rect 182639 290869 182667 290897
rect 182701 290869 182729 290897
rect 182763 290869 182791 290897
rect 182577 290807 182605 290835
rect 182639 290807 182667 290835
rect 182701 290807 182729 290835
rect 182763 290807 182791 290835
rect 182577 290745 182605 290773
rect 182639 290745 182667 290773
rect 182701 290745 182729 290773
rect 182763 290745 182791 290773
rect 182577 281931 182605 281959
rect 182639 281931 182667 281959
rect 182701 281931 182729 281959
rect 182763 281931 182791 281959
rect 182577 281869 182605 281897
rect 182639 281869 182667 281897
rect 182701 281869 182729 281897
rect 182763 281869 182791 281897
rect 182577 281807 182605 281835
rect 182639 281807 182667 281835
rect 182701 281807 182729 281835
rect 182763 281807 182791 281835
rect 182577 281745 182605 281773
rect 182639 281745 182667 281773
rect 182701 281745 182729 281773
rect 182763 281745 182791 281773
rect 182577 272931 182605 272959
rect 182639 272931 182667 272959
rect 182701 272931 182729 272959
rect 182763 272931 182791 272959
rect 182577 272869 182605 272897
rect 182639 272869 182667 272897
rect 182701 272869 182729 272897
rect 182763 272869 182791 272897
rect 182577 272807 182605 272835
rect 182639 272807 182667 272835
rect 182701 272807 182729 272835
rect 182763 272807 182791 272835
rect 182577 272745 182605 272773
rect 182639 272745 182667 272773
rect 182701 272745 182729 272773
rect 182763 272745 182791 272773
rect 182577 263931 182605 263959
rect 182639 263931 182667 263959
rect 182701 263931 182729 263959
rect 182763 263931 182791 263959
rect 182577 263869 182605 263897
rect 182639 263869 182667 263897
rect 182701 263869 182729 263897
rect 182763 263869 182791 263897
rect 182577 263807 182605 263835
rect 182639 263807 182667 263835
rect 182701 263807 182729 263835
rect 182763 263807 182791 263835
rect 182577 263745 182605 263773
rect 182639 263745 182667 263773
rect 182701 263745 182729 263773
rect 182763 263745 182791 263773
rect 182577 254931 182605 254959
rect 182639 254931 182667 254959
rect 182701 254931 182729 254959
rect 182763 254931 182791 254959
rect 182577 254869 182605 254897
rect 182639 254869 182667 254897
rect 182701 254869 182729 254897
rect 182763 254869 182791 254897
rect 182577 254807 182605 254835
rect 182639 254807 182667 254835
rect 182701 254807 182729 254835
rect 182763 254807 182791 254835
rect 182577 254745 182605 254773
rect 182639 254745 182667 254773
rect 182701 254745 182729 254773
rect 182763 254745 182791 254773
rect 184437 299642 184465 299670
rect 184499 299642 184527 299670
rect 184561 299642 184589 299670
rect 184623 299642 184651 299670
rect 184437 299580 184465 299608
rect 184499 299580 184527 299608
rect 184561 299580 184589 299608
rect 184623 299580 184651 299608
rect 184437 299518 184465 299546
rect 184499 299518 184527 299546
rect 184561 299518 184589 299546
rect 184623 299518 184651 299546
rect 184437 299456 184465 299484
rect 184499 299456 184527 299484
rect 184561 299456 184589 299484
rect 184623 299456 184651 299484
rect 184437 293931 184465 293959
rect 184499 293931 184527 293959
rect 184561 293931 184589 293959
rect 184623 293931 184651 293959
rect 184437 293869 184465 293897
rect 184499 293869 184527 293897
rect 184561 293869 184589 293897
rect 184623 293869 184651 293897
rect 184437 293807 184465 293835
rect 184499 293807 184527 293835
rect 184561 293807 184589 293835
rect 184623 293807 184651 293835
rect 184437 293745 184465 293773
rect 184499 293745 184527 293773
rect 184561 293745 184589 293773
rect 184623 293745 184651 293773
rect 184437 284931 184465 284959
rect 184499 284931 184527 284959
rect 184561 284931 184589 284959
rect 184623 284931 184651 284959
rect 184437 284869 184465 284897
rect 184499 284869 184527 284897
rect 184561 284869 184589 284897
rect 184623 284869 184651 284897
rect 184437 284807 184465 284835
rect 184499 284807 184527 284835
rect 184561 284807 184589 284835
rect 184623 284807 184651 284835
rect 184437 284745 184465 284773
rect 184499 284745 184527 284773
rect 184561 284745 184589 284773
rect 184623 284745 184651 284773
rect 184437 275931 184465 275959
rect 184499 275931 184527 275959
rect 184561 275931 184589 275959
rect 184623 275931 184651 275959
rect 184437 275869 184465 275897
rect 184499 275869 184527 275897
rect 184561 275869 184589 275897
rect 184623 275869 184651 275897
rect 184437 275807 184465 275835
rect 184499 275807 184527 275835
rect 184561 275807 184589 275835
rect 184623 275807 184651 275835
rect 184437 275745 184465 275773
rect 184499 275745 184527 275773
rect 184561 275745 184589 275773
rect 184623 275745 184651 275773
rect 184437 266931 184465 266959
rect 184499 266931 184527 266959
rect 184561 266931 184589 266959
rect 184623 266931 184651 266959
rect 184437 266869 184465 266897
rect 184499 266869 184527 266897
rect 184561 266869 184589 266897
rect 184623 266869 184651 266897
rect 184437 266807 184465 266835
rect 184499 266807 184527 266835
rect 184561 266807 184589 266835
rect 184623 266807 184651 266835
rect 184437 266745 184465 266773
rect 184499 266745 184527 266773
rect 184561 266745 184589 266773
rect 184623 266745 184651 266773
rect 184437 257931 184465 257959
rect 184499 257931 184527 257959
rect 184561 257931 184589 257959
rect 184623 257931 184651 257959
rect 184437 257869 184465 257897
rect 184499 257869 184527 257897
rect 184561 257869 184589 257897
rect 184623 257869 184651 257897
rect 184437 257807 184465 257835
rect 184499 257807 184527 257835
rect 184561 257807 184589 257835
rect 184623 257807 184651 257835
rect 184437 257745 184465 257773
rect 184499 257745 184527 257773
rect 184561 257745 184589 257773
rect 184623 257745 184651 257773
rect 191577 299162 191605 299190
rect 191639 299162 191667 299190
rect 191701 299162 191729 299190
rect 191763 299162 191791 299190
rect 191577 299100 191605 299128
rect 191639 299100 191667 299128
rect 191701 299100 191729 299128
rect 191763 299100 191791 299128
rect 191577 299038 191605 299066
rect 191639 299038 191667 299066
rect 191701 299038 191729 299066
rect 191763 299038 191791 299066
rect 191577 298976 191605 299004
rect 191639 298976 191667 299004
rect 191701 298976 191729 299004
rect 191763 298976 191791 299004
rect 191577 290931 191605 290959
rect 191639 290931 191667 290959
rect 191701 290931 191729 290959
rect 191763 290931 191791 290959
rect 191577 290869 191605 290897
rect 191639 290869 191667 290897
rect 191701 290869 191729 290897
rect 191763 290869 191791 290897
rect 191577 290807 191605 290835
rect 191639 290807 191667 290835
rect 191701 290807 191729 290835
rect 191763 290807 191791 290835
rect 191577 290745 191605 290773
rect 191639 290745 191667 290773
rect 191701 290745 191729 290773
rect 191763 290745 191791 290773
rect 191577 281931 191605 281959
rect 191639 281931 191667 281959
rect 191701 281931 191729 281959
rect 191763 281931 191791 281959
rect 191577 281869 191605 281897
rect 191639 281869 191667 281897
rect 191701 281869 191729 281897
rect 191763 281869 191791 281897
rect 191577 281807 191605 281835
rect 191639 281807 191667 281835
rect 191701 281807 191729 281835
rect 191763 281807 191791 281835
rect 191577 281745 191605 281773
rect 191639 281745 191667 281773
rect 191701 281745 191729 281773
rect 191763 281745 191791 281773
rect 191577 272931 191605 272959
rect 191639 272931 191667 272959
rect 191701 272931 191729 272959
rect 191763 272931 191791 272959
rect 191577 272869 191605 272897
rect 191639 272869 191667 272897
rect 191701 272869 191729 272897
rect 191763 272869 191791 272897
rect 191577 272807 191605 272835
rect 191639 272807 191667 272835
rect 191701 272807 191729 272835
rect 191763 272807 191791 272835
rect 191577 272745 191605 272773
rect 191639 272745 191667 272773
rect 191701 272745 191729 272773
rect 191763 272745 191791 272773
rect 191577 263931 191605 263959
rect 191639 263931 191667 263959
rect 191701 263931 191729 263959
rect 191763 263931 191791 263959
rect 191577 263869 191605 263897
rect 191639 263869 191667 263897
rect 191701 263869 191729 263897
rect 191763 263869 191791 263897
rect 191577 263807 191605 263835
rect 191639 263807 191667 263835
rect 191701 263807 191729 263835
rect 191763 263807 191791 263835
rect 191577 263745 191605 263773
rect 191639 263745 191667 263773
rect 191701 263745 191729 263773
rect 191763 263745 191791 263773
rect 191577 254931 191605 254959
rect 191639 254931 191667 254959
rect 191701 254931 191729 254959
rect 191763 254931 191791 254959
rect 191577 254869 191605 254897
rect 191639 254869 191667 254897
rect 191701 254869 191729 254897
rect 191763 254869 191791 254897
rect 191577 254807 191605 254835
rect 191639 254807 191667 254835
rect 191701 254807 191729 254835
rect 191763 254807 191791 254835
rect 191577 254745 191605 254773
rect 191639 254745 191667 254773
rect 191701 254745 191729 254773
rect 191763 254745 191791 254773
rect 193437 299642 193465 299670
rect 193499 299642 193527 299670
rect 193561 299642 193589 299670
rect 193623 299642 193651 299670
rect 193437 299580 193465 299608
rect 193499 299580 193527 299608
rect 193561 299580 193589 299608
rect 193623 299580 193651 299608
rect 193437 299518 193465 299546
rect 193499 299518 193527 299546
rect 193561 299518 193589 299546
rect 193623 299518 193651 299546
rect 193437 299456 193465 299484
rect 193499 299456 193527 299484
rect 193561 299456 193589 299484
rect 193623 299456 193651 299484
rect 193437 293931 193465 293959
rect 193499 293931 193527 293959
rect 193561 293931 193589 293959
rect 193623 293931 193651 293959
rect 193437 293869 193465 293897
rect 193499 293869 193527 293897
rect 193561 293869 193589 293897
rect 193623 293869 193651 293897
rect 193437 293807 193465 293835
rect 193499 293807 193527 293835
rect 193561 293807 193589 293835
rect 193623 293807 193651 293835
rect 193437 293745 193465 293773
rect 193499 293745 193527 293773
rect 193561 293745 193589 293773
rect 193623 293745 193651 293773
rect 193437 284931 193465 284959
rect 193499 284931 193527 284959
rect 193561 284931 193589 284959
rect 193623 284931 193651 284959
rect 193437 284869 193465 284897
rect 193499 284869 193527 284897
rect 193561 284869 193589 284897
rect 193623 284869 193651 284897
rect 193437 284807 193465 284835
rect 193499 284807 193527 284835
rect 193561 284807 193589 284835
rect 193623 284807 193651 284835
rect 193437 284745 193465 284773
rect 193499 284745 193527 284773
rect 193561 284745 193589 284773
rect 193623 284745 193651 284773
rect 193437 275931 193465 275959
rect 193499 275931 193527 275959
rect 193561 275931 193589 275959
rect 193623 275931 193651 275959
rect 193437 275869 193465 275897
rect 193499 275869 193527 275897
rect 193561 275869 193589 275897
rect 193623 275869 193651 275897
rect 193437 275807 193465 275835
rect 193499 275807 193527 275835
rect 193561 275807 193589 275835
rect 193623 275807 193651 275835
rect 193437 275745 193465 275773
rect 193499 275745 193527 275773
rect 193561 275745 193589 275773
rect 193623 275745 193651 275773
rect 193437 266931 193465 266959
rect 193499 266931 193527 266959
rect 193561 266931 193589 266959
rect 193623 266931 193651 266959
rect 193437 266869 193465 266897
rect 193499 266869 193527 266897
rect 193561 266869 193589 266897
rect 193623 266869 193651 266897
rect 193437 266807 193465 266835
rect 193499 266807 193527 266835
rect 193561 266807 193589 266835
rect 193623 266807 193651 266835
rect 193437 266745 193465 266773
rect 193499 266745 193527 266773
rect 193561 266745 193589 266773
rect 193623 266745 193651 266773
rect 193437 257931 193465 257959
rect 193499 257931 193527 257959
rect 193561 257931 193589 257959
rect 193623 257931 193651 257959
rect 193437 257869 193465 257897
rect 193499 257869 193527 257897
rect 193561 257869 193589 257897
rect 193623 257869 193651 257897
rect 193437 257807 193465 257835
rect 193499 257807 193527 257835
rect 193561 257807 193589 257835
rect 193623 257807 193651 257835
rect 193437 257745 193465 257773
rect 193499 257745 193527 257773
rect 193561 257745 193589 257773
rect 193623 257745 193651 257773
rect 200577 299162 200605 299190
rect 200639 299162 200667 299190
rect 200701 299162 200729 299190
rect 200763 299162 200791 299190
rect 200577 299100 200605 299128
rect 200639 299100 200667 299128
rect 200701 299100 200729 299128
rect 200763 299100 200791 299128
rect 200577 299038 200605 299066
rect 200639 299038 200667 299066
rect 200701 299038 200729 299066
rect 200763 299038 200791 299066
rect 200577 298976 200605 299004
rect 200639 298976 200667 299004
rect 200701 298976 200729 299004
rect 200763 298976 200791 299004
rect 200577 290931 200605 290959
rect 200639 290931 200667 290959
rect 200701 290931 200729 290959
rect 200763 290931 200791 290959
rect 200577 290869 200605 290897
rect 200639 290869 200667 290897
rect 200701 290869 200729 290897
rect 200763 290869 200791 290897
rect 200577 290807 200605 290835
rect 200639 290807 200667 290835
rect 200701 290807 200729 290835
rect 200763 290807 200791 290835
rect 200577 290745 200605 290773
rect 200639 290745 200667 290773
rect 200701 290745 200729 290773
rect 200763 290745 200791 290773
rect 200577 281931 200605 281959
rect 200639 281931 200667 281959
rect 200701 281931 200729 281959
rect 200763 281931 200791 281959
rect 200577 281869 200605 281897
rect 200639 281869 200667 281897
rect 200701 281869 200729 281897
rect 200763 281869 200791 281897
rect 200577 281807 200605 281835
rect 200639 281807 200667 281835
rect 200701 281807 200729 281835
rect 200763 281807 200791 281835
rect 200577 281745 200605 281773
rect 200639 281745 200667 281773
rect 200701 281745 200729 281773
rect 200763 281745 200791 281773
rect 200577 272931 200605 272959
rect 200639 272931 200667 272959
rect 200701 272931 200729 272959
rect 200763 272931 200791 272959
rect 200577 272869 200605 272897
rect 200639 272869 200667 272897
rect 200701 272869 200729 272897
rect 200763 272869 200791 272897
rect 200577 272807 200605 272835
rect 200639 272807 200667 272835
rect 200701 272807 200729 272835
rect 200763 272807 200791 272835
rect 200577 272745 200605 272773
rect 200639 272745 200667 272773
rect 200701 272745 200729 272773
rect 200763 272745 200791 272773
rect 200577 263931 200605 263959
rect 200639 263931 200667 263959
rect 200701 263931 200729 263959
rect 200763 263931 200791 263959
rect 200577 263869 200605 263897
rect 200639 263869 200667 263897
rect 200701 263869 200729 263897
rect 200763 263869 200791 263897
rect 200577 263807 200605 263835
rect 200639 263807 200667 263835
rect 200701 263807 200729 263835
rect 200763 263807 200791 263835
rect 200577 263745 200605 263773
rect 200639 263745 200667 263773
rect 200701 263745 200729 263773
rect 200763 263745 200791 263773
rect 200577 254931 200605 254959
rect 200639 254931 200667 254959
rect 200701 254931 200729 254959
rect 200763 254931 200791 254959
rect 200577 254869 200605 254897
rect 200639 254869 200667 254897
rect 200701 254869 200729 254897
rect 200763 254869 200791 254897
rect 200577 254807 200605 254835
rect 200639 254807 200667 254835
rect 200701 254807 200729 254835
rect 200763 254807 200791 254835
rect 200577 254745 200605 254773
rect 200639 254745 200667 254773
rect 200701 254745 200729 254773
rect 200763 254745 200791 254773
rect 202437 299642 202465 299670
rect 202499 299642 202527 299670
rect 202561 299642 202589 299670
rect 202623 299642 202651 299670
rect 202437 299580 202465 299608
rect 202499 299580 202527 299608
rect 202561 299580 202589 299608
rect 202623 299580 202651 299608
rect 202437 299518 202465 299546
rect 202499 299518 202527 299546
rect 202561 299518 202589 299546
rect 202623 299518 202651 299546
rect 202437 299456 202465 299484
rect 202499 299456 202527 299484
rect 202561 299456 202589 299484
rect 202623 299456 202651 299484
rect 202437 293931 202465 293959
rect 202499 293931 202527 293959
rect 202561 293931 202589 293959
rect 202623 293931 202651 293959
rect 202437 293869 202465 293897
rect 202499 293869 202527 293897
rect 202561 293869 202589 293897
rect 202623 293869 202651 293897
rect 202437 293807 202465 293835
rect 202499 293807 202527 293835
rect 202561 293807 202589 293835
rect 202623 293807 202651 293835
rect 202437 293745 202465 293773
rect 202499 293745 202527 293773
rect 202561 293745 202589 293773
rect 202623 293745 202651 293773
rect 202437 284931 202465 284959
rect 202499 284931 202527 284959
rect 202561 284931 202589 284959
rect 202623 284931 202651 284959
rect 202437 284869 202465 284897
rect 202499 284869 202527 284897
rect 202561 284869 202589 284897
rect 202623 284869 202651 284897
rect 202437 284807 202465 284835
rect 202499 284807 202527 284835
rect 202561 284807 202589 284835
rect 202623 284807 202651 284835
rect 202437 284745 202465 284773
rect 202499 284745 202527 284773
rect 202561 284745 202589 284773
rect 202623 284745 202651 284773
rect 202437 275931 202465 275959
rect 202499 275931 202527 275959
rect 202561 275931 202589 275959
rect 202623 275931 202651 275959
rect 202437 275869 202465 275897
rect 202499 275869 202527 275897
rect 202561 275869 202589 275897
rect 202623 275869 202651 275897
rect 202437 275807 202465 275835
rect 202499 275807 202527 275835
rect 202561 275807 202589 275835
rect 202623 275807 202651 275835
rect 202437 275745 202465 275773
rect 202499 275745 202527 275773
rect 202561 275745 202589 275773
rect 202623 275745 202651 275773
rect 202437 266931 202465 266959
rect 202499 266931 202527 266959
rect 202561 266931 202589 266959
rect 202623 266931 202651 266959
rect 202437 266869 202465 266897
rect 202499 266869 202527 266897
rect 202561 266869 202589 266897
rect 202623 266869 202651 266897
rect 202437 266807 202465 266835
rect 202499 266807 202527 266835
rect 202561 266807 202589 266835
rect 202623 266807 202651 266835
rect 202437 266745 202465 266773
rect 202499 266745 202527 266773
rect 202561 266745 202589 266773
rect 202623 266745 202651 266773
rect 202437 257931 202465 257959
rect 202499 257931 202527 257959
rect 202561 257931 202589 257959
rect 202623 257931 202651 257959
rect 202437 257869 202465 257897
rect 202499 257869 202527 257897
rect 202561 257869 202589 257897
rect 202623 257869 202651 257897
rect 202437 257807 202465 257835
rect 202499 257807 202527 257835
rect 202561 257807 202589 257835
rect 202623 257807 202651 257835
rect 202437 257745 202465 257773
rect 202499 257745 202527 257773
rect 202561 257745 202589 257773
rect 202623 257745 202651 257773
rect 209577 299162 209605 299190
rect 209639 299162 209667 299190
rect 209701 299162 209729 299190
rect 209763 299162 209791 299190
rect 209577 299100 209605 299128
rect 209639 299100 209667 299128
rect 209701 299100 209729 299128
rect 209763 299100 209791 299128
rect 209577 299038 209605 299066
rect 209639 299038 209667 299066
rect 209701 299038 209729 299066
rect 209763 299038 209791 299066
rect 209577 298976 209605 299004
rect 209639 298976 209667 299004
rect 209701 298976 209729 299004
rect 209763 298976 209791 299004
rect 209577 290931 209605 290959
rect 209639 290931 209667 290959
rect 209701 290931 209729 290959
rect 209763 290931 209791 290959
rect 209577 290869 209605 290897
rect 209639 290869 209667 290897
rect 209701 290869 209729 290897
rect 209763 290869 209791 290897
rect 209577 290807 209605 290835
rect 209639 290807 209667 290835
rect 209701 290807 209729 290835
rect 209763 290807 209791 290835
rect 209577 290745 209605 290773
rect 209639 290745 209667 290773
rect 209701 290745 209729 290773
rect 209763 290745 209791 290773
rect 209577 281931 209605 281959
rect 209639 281931 209667 281959
rect 209701 281931 209729 281959
rect 209763 281931 209791 281959
rect 209577 281869 209605 281897
rect 209639 281869 209667 281897
rect 209701 281869 209729 281897
rect 209763 281869 209791 281897
rect 209577 281807 209605 281835
rect 209639 281807 209667 281835
rect 209701 281807 209729 281835
rect 209763 281807 209791 281835
rect 209577 281745 209605 281773
rect 209639 281745 209667 281773
rect 209701 281745 209729 281773
rect 209763 281745 209791 281773
rect 209577 272931 209605 272959
rect 209639 272931 209667 272959
rect 209701 272931 209729 272959
rect 209763 272931 209791 272959
rect 209577 272869 209605 272897
rect 209639 272869 209667 272897
rect 209701 272869 209729 272897
rect 209763 272869 209791 272897
rect 209577 272807 209605 272835
rect 209639 272807 209667 272835
rect 209701 272807 209729 272835
rect 209763 272807 209791 272835
rect 209577 272745 209605 272773
rect 209639 272745 209667 272773
rect 209701 272745 209729 272773
rect 209763 272745 209791 272773
rect 209577 263931 209605 263959
rect 209639 263931 209667 263959
rect 209701 263931 209729 263959
rect 209763 263931 209791 263959
rect 209577 263869 209605 263897
rect 209639 263869 209667 263897
rect 209701 263869 209729 263897
rect 209763 263869 209791 263897
rect 209577 263807 209605 263835
rect 209639 263807 209667 263835
rect 209701 263807 209729 263835
rect 209763 263807 209791 263835
rect 209577 263745 209605 263773
rect 209639 263745 209667 263773
rect 209701 263745 209729 263773
rect 209763 263745 209791 263773
rect 209577 254931 209605 254959
rect 209639 254931 209667 254959
rect 209701 254931 209729 254959
rect 209763 254931 209791 254959
rect 209577 254869 209605 254897
rect 209639 254869 209667 254897
rect 209701 254869 209729 254897
rect 209763 254869 209791 254897
rect 209577 254807 209605 254835
rect 209639 254807 209667 254835
rect 209701 254807 209729 254835
rect 209763 254807 209791 254835
rect 209577 254745 209605 254773
rect 209639 254745 209667 254773
rect 209701 254745 209729 254773
rect 209763 254745 209791 254773
rect 211437 299642 211465 299670
rect 211499 299642 211527 299670
rect 211561 299642 211589 299670
rect 211623 299642 211651 299670
rect 211437 299580 211465 299608
rect 211499 299580 211527 299608
rect 211561 299580 211589 299608
rect 211623 299580 211651 299608
rect 211437 299518 211465 299546
rect 211499 299518 211527 299546
rect 211561 299518 211589 299546
rect 211623 299518 211651 299546
rect 211437 299456 211465 299484
rect 211499 299456 211527 299484
rect 211561 299456 211589 299484
rect 211623 299456 211651 299484
rect 211437 293931 211465 293959
rect 211499 293931 211527 293959
rect 211561 293931 211589 293959
rect 211623 293931 211651 293959
rect 211437 293869 211465 293897
rect 211499 293869 211527 293897
rect 211561 293869 211589 293897
rect 211623 293869 211651 293897
rect 211437 293807 211465 293835
rect 211499 293807 211527 293835
rect 211561 293807 211589 293835
rect 211623 293807 211651 293835
rect 211437 293745 211465 293773
rect 211499 293745 211527 293773
rect 211561 293745 211589 293773
rect 211623 293745 211651 293773
rect 211437 284931 211465 284959
rect 211499 284931 211527 284959
rect 211561 284931 211589 284959
rect 211623 284931 211651 284959
rect 211437 284869 211465 284897
rect 211499 284869 211527 284897
rect 211561 284869 211589 284897
rect 211623 284869 211651 284897
rect 211437 284807 211465 284835
rect 211499 284807 211527 284835
rect 211561 284807 211589 284835
rect 211623 284807 211651 284835
rect 211437 284745 211465 284773
rect 211499 284745 211527 284773
rect 211561 284745 211589 284773
rect 211623 284745 211651 284773
rect 211437 275931 211465 275959
rect 211499 275931 211527 275959
rect 211561 275931 211589 275959
rect 211623 275931 211651 275959
rect 211437 275869 211465 275897
rect 211499 275869 211527 275897
rect 211561 275869 211589 275897
rect 211623 275869 211651 275897
rect 211437 275807 211465 275835
rect 211499 275807 211527 275835
rect 211561 275807 211589 275835
rect 211623 275807 211651 275835
rect 211437 275745 211465 275773
rect 211499 275745 211527 275773
rect 211561 275745 211589 275773
rect 211623 275745 211651 275773
rect 211437 266931 211465 266959
rect 211499 266931 211527 266959
rect 211561 266931 211589 266959
rect 211623 266931 211651 266959
rect 211437 266869 211465 266897
rect 211499 266869 211527 266897
rect 211561 266869 211589 266897
rect 211623 266869 211651 266897
rect 211437 266807 211465 266835
rect 211499 266807 211527 266835
rect 211561 266807 211589 266835
rect 211623 266807 211651 266835
rect 211437 266745 211465 266773
rect 211499 266745 211527 266773
rect 211561 266745 211589 266773
rect 211623 266745 211651 266773
rect 211437 257931 211465 257959
rect 211499 257931 211527 257959
rect 211561 257931 211589 257959
rect 211623 257931 211651 257959
rect 211437 257869 211465 257897
rect 211499 257869 211527 257897
rect 211561 257869 211589 257897
rect 211623 257869 211651 257897
rect 211437 257807 211465 257835
rect 211499 257807 211527 257835
rect 211561 257807 211589 257835
rect 211623 257807 211651 257835
rect 211437 257745 211465 257773
rect 211499 257745 211527 257773
rect 211561 257745 211589 257773
rect 211623 257745 211651 257773
rect 218577 299162 218605 299190
rect 218639 299162 218667 299190
rect 218701 299162 218729 299190
rect 218763 299162 218791 299190
rect 218577 299100 218605 299128
rect 218639 299100 218667 299128
rect 218701 299100 218729 299128
rect 218763 299100 218791 299128
rect 218577 299038 218605 299066
rect 218639 299038 218667 299066
rect 218701 299038 218729 299066
rect 218763 299038 218791 299066
rect 218577 298976 218605 299004
rect 218639 298976 218667 299004
rect 218701 298976 218729 299004
rect 218763 298976 218791 299004
rect 218577 290931 218605 290959
rect 218639 290931 218667 290959
rect 218701 290931 218729 290959
rect 218763 290931 218791 290959
rect 218577 290869 218605 290897
rect 218639 290869 218667 290897
rect 218701 290869 218729 290897
rect 218763 290869 218791 290897
rect 218577 290807 218605 290835
rect 218639 290807 218667 290835
rect 218701 290807 218729 290835
rect 218763 290807 218791 290835
rect 218577 290745 218605 290773
rect 218639 290745 218667 290773
rect 218701 290745 218729 290773
rect 218763 290745 218791 290773
rect 218577 281931 218605 281959
rect 218639 281931 218667 281959
rect 218701 281931 218729 281959
rect 218763 281931 218791 281959
rect 218577 281869 218605 281897
rect 218639 281869 218667 281897
rect 218701 281869 218729 281897
rect 218763 281869 218791 281897
rect 218577 281807 218605 281835
rect 218639 281807 218667 281835
rect 218701 281807 218729 281835
rect 218763 281807 218791 281835
rect 218577 281745 218605 281773
rect 218639 281745 218667 281773
rect 218701 281745 218729 281773
rect 218763 281745 218791 281773
rect 218577 272931 218605 272959
rect 218639 272931 218667 272959
rect 218701 272931 218729 272959
rect 218763 272931 218791 272959
rect 218577 272869 218605 272897
rect 218639 272869 218667 272897
rect 218701 272869 218729 272897
rect 218763 272869 218791 272897
rect 218577 272807 218605 272835
rect 218639 272807 218667 272835
rect 218701 272807 218729 272835
rect 218763 272807 218791 272835
rect 218577 272745 218605 272773
rect 218639 272745 218667 272773
rect 218701 272745 218729 272773
rect 218763 272745 218791 272773
rect 218577 263931 218605 263959
rect 218639 263931 218667 263959
rect 218701 263931 218729 263959
rect 218763 263931 218791 263959
rect 218577 263869 218605 263897
rect 218639 263869 218667 263897
rect 218701 263869 218729 263897
rect 218763 263869 218791 263897
rect 218577 263807 218605 263835
rect 218639 263807 218667 263835
rect 218701 263807 218729 263835
rect 218763 263807 218791 263835
rect 218577 263745 218605 263773
rect 218639 263745 218667 263773
rect 218701 263745 218729 263773
rect 218763 263745 218791 263773
rect 218577 254931 218605 254959
rect 218639 254931 218667 254959
rect 218701 254931 218729 254959
rect 218763 254931 218791 254959
rect 218577 254869 218605 254897
rect 218639 254869 218667 254897
rect 218701 254869 218729 254897
rect 218763 254869 218791 254897
rect 218577 254807 218605 254835
rect 218639 254807 218667 254835
rect 218701 254807 218729 254835
rect 218763 254807 218791 254835
rect 218577 254745 218605 254773
rect 218639 254745 218667 254773
rect 218701 254745 218729 254773
rect 218763 254745 218791 254773
rect 220437 299642 220465 299670
rect 220499 299642 220527 299670
rect 220561 299642 220589 299670
rect 220623 299642 220651 299670
rect 220437 299580 220465 299608
rect 220499 299580 220527 299608
rect 220561 299580 220589 299608
rect 220623 299580 220651 299608
rect 220437 299518 220465 299546
rect 220499 299518 220527 299546
rect 220561 299518 220589 299546
rect 220623 299518 220651 299546
rect 220437 299456 220465 299484
rect 220499 299456 220527 299484
rect 220561 299456 220589 299484
rect 220623 299456 220651 299484
rect 220437 293931 220465 293959
rect 220499 293931 220527 293959
rect 220561 293931 220589 293959
rect 220623 293931 220651 293959
rect 220437 293869 220465 293897
rect 220499 293869 220527 293897
rect 220561 293869 220589 293897
rect 220623 293869 220651 293897
rect 220437 293807 220465 293835
rect 220499 293807 220527 293835
rect 220561 293807 220589 293835
rect 220623 293807 220651 293835
rect 220437 293745 220465 293773
rect 220499 293745 220527 293773
rect 220561 293745 220589 293773
rect 220623 293745 220651 293773
rect 220437 284931 220465 284959
rect 220499 284931 220527 284959
rect 220561 284931 220589 284959
rect 220623 284931 220651 284959
rect 220437 284869 220465 284897
rect 220499 284869 220527 284897
rect 220561 284869 220589 284897
rect 220623 284869 220651 284897
rect 220437 284807 220465 284835
rect 220499 284807 220527 284835
rect 220561 284807 220589 284835
rect 220623 284807 220651 284835
rect 220437 284745 220465 284773
rect 220499 284745 220527 284773
rect 220561 284745 220589 284773
rect 220623 284745 220651 284773
rect 220437 275931 220465 275959
rect 220499 275931 220527 275959
rect 220561 275931 220589 275959
rect 220623 275931 220651 275959
rect 220437 275869 220465 275897
rect 220499 275869 220527 275897
rect 220561 275869 220589 275897
rect 220623 275869 220651 275897
rect 220437 275807 220465 275835
rect 220499 275807 220527 275835
rect 220561 275807 220589 275835
rect 220623 275807 220651 275835
rect 220437 275745 220465 275773
rect 220499 275745 220527 275773
rect 220561 275745 220589 275773
rect 220623 275745 220651 275773
rect 220437 266931 220465 266959
rect 220499 266931 220527 266959
rect 220561 266931 220589 266959
rect 220623 266931 220651 266959
rect 220437 266869 220465 266897
rect 220499 266869 220527 266897
rect 220561 266869 220589 266897
rect 220623 266869 220651 266897
rect 220437 266807 220465 266835
rect 220499 266807 220527 266835
rect 220561 266807 220589 266835
rect 220623 266807 220651 266835
rect 220437 266745 220465 266773
rect 220499 266745 220527 266773
rect 220561 266745 220589 266773
rect 220623 266745 220651 266773
rect 220437 257931 220465 257959
rect 220499 257931 220527 257959
rect 220561 257931 220589 257959
rect 220623 257931 220651 257959
rect 220437 257869 220465 257897
rect 220499 257869 220527 257897
rect 220561 257869 220589 257897
rect 220623 257869 220651 257897
rect 220437 257807 220465 257835
rect 220499 257807 220527 257835
rect 220561 257807 220589 257835
rect 220623 257807 220651 257835
rect 220437 257745 220465 257773
rect 220499 257745 220527 257773
rect 220561 257745 220589 257773
rect 220623 257745 220651 257773
rect 227577 299162 227605 299190
rect 227639 299162 227667 299190
rect 227701 299162 227729 299190
rect 227763 299162 227791 299190
rect 227577 299100 227605 299128
rect 227639 299100 227667 299128
rect 227701 299100 227729 299128
rect 227763 299100 227791 299128
rect 227577 299038 227605 299066
rect 227639 299038 227667 299066
rect 227701 299038 227729 299066
rect 227763 299038 227791 299066
rect 227577 298976 227605 299004
rect 227639 298976 227667 299004
rect 227701 298976 227729 299004
rect 227763 298976 227791 299004
rect 227577 290931 227605 290959
rect 227639 290931 227667 290959
rect 227701 290931 227729 290959
rect 227763 290931 227791 290959
rect 227577 290869 227605 290897
rect 227639 290869 227667 290897
rect 227701 290869 227729 290897
rect 227763 290869 227791 290897
rect 227577 290807 227605 290835
rect 227639 290807 227667 290835
rect 227701 290807 227729 290835
rect 227763 290807 227791 290835
rect 227577 290745 227605 290773
rect 227639 290745 227667 290773
rect 227701 290745 227729 290773
rect 227763 290745 227791 290773
rect 227577 281931 227605 281959
rect 227639 281931 227667 281959
rect 227701 281931 227729 281959
rect 227763 281931 227791 281959
rect 227577 281869 227605 281897
rect 227639 281869 227667 281897
rect 227701 281869 227729 281897
rect 227763 281869 227791 281897
rect 227577 281807 227605 281835
rect 227639 281807 227667 281835
rect 227701 281807 227729 281835
rect 227763 281807 227791 281835
rect 227577 281745 227605 281773
rect 227639 281745 227667 281773
rect 227701 281745 227729 281773
rect 227763 281745 227791 281773
rect 227577 272931 227605 272959
rect 227639 272931 227667 272959
rect 227701 272931 227729 272959
rect 227763 272931 227791 272959
rect 227577 272869 227605 272897
rect 227639 272869 227667 272897
rect 227701 272869 227729 272897
rect 227763 272869 227791 272897
rect 227577 272807 227605 272835
rect 227639 272807 227667 272835
rect 227701 272807 227729 272835
rect 227763 272807 227791 272835
rect 227577 272745 227605 272773
rect 227639 272745 227667 272773
rect 227701 272745 227729 272773
rect 227763 272745 227791 272773
rect 227577 263931 227605 263959
rect 227639 263931 227667 263959
rect 227701 263931 227729 263959
rect 227763 263931 227791 263959
rect 227577 263869 227605 263897
rect 227639 263869 227667 263897
rect 227701 263869 227729 263897
rect 227763 263869 227791 263897
rect 227577 263807 227605 263835
rect 227639 263807 227667 263835
rect 227701 263807 227729 263835
rect 227763 263807 227791 263835
rect 227577 263745 227605 263773
rect 227639 263745 227667 263773
rect 227701 263745 227729 263773
rect 227763 263745 227791 263773
rect 227577 254931 227605 254959
rect 227639 254931 227667 254959
rect 227701 254931 227729 254959
rect 227763 254931 227791 254959
rect 227577 254869 227605 254897
rect 227639 254869 227667 254897
rect 227701 254869 227729 254897
rect 227763 254869 227791 254897
rect 227577 254807 227605 254835
rect 227639 254807 227667 254835
rect 227701 254807 227729 254835
rect 227763 254807 227791 254835
rect 227577 254745 227605 254773
rect 227639 254745 227667 254773
rect 227701 254745 227729 254773
rect 227763 254745 227791 254773
rect 229437 299642 229465 299670
rect 229499 299642 229527 299670
rect 229561 299642 229589 299670
rect 229623 299642 229651 299670
rect 229437 299580 229465 299608
rect 229499 299580 229527 299608
rect 229561 299580 229589 299608
rect 229623 299580 229651 299608
rect 229437 299518 229465 299546
rect 229499 299518 229527 299546
rect 229561 299518 229589 299546
rect 229623 299518 229651 299546
rect 229437 299456 229465 299484
rect 229499 299456 229527 299484
rect 229561 299456 229589 299484
rect 229623 299456 229651 299484
rect 229437 293931 229465 293959
rect 229499 293931 229527 293959
rect 229561 293931 229589 293959
rect 229623 293931 229651 293959
rect 229437 293869 229465 293897
rect 229499 293869 229527 293897
rect 229561 293869 229589 293897
rect 229623 293869 229651 293897
rect 229437 293807 229465 293835
rect 229499 293807 229527 293835
rect 229561 293807 229589 293835
rect 229623 293807 229651 293835
rect 229437 293745 229465 293773
rect 229499 293745 229527 293773
rect 229561 293745 229589 293773
rect 229623 293745 229651 293773
rect 229437 284931 229465 284959
rect 229499 284931 229527 284959
rect 229561 284931 229589 284959
rect 229623 284931 229651 284959
rect 229437 284869 229465 284897
rect 229499 284869 229527 284897
rect 229561 284869 229589 284897
rect 229623 284869 229651 284897
rect 229437 284807 229465 284835
rect 229499 284807 229527 284835
rect 229561 284807 229589 284835
rect 229623 284807 229651 284835
rect 229437 284745 229465 284773
rect 229499 284745 229527 284773
rect 229561 284745 229589 284773
rect 229623 284745 229651 284773
rect 229437 275931 229465 275959
rect 229499 275931 229527 275959
rect 229561 275931 229589 275959
rect 229623 275931 229651 275959
rect 229437 275869 229465 275897
rect 229499 275869 229527 275897
rect 229561 275869 229589 275897
rect 229623 275869 229651 275897
rect 229437 275807 229465 275835
rect 229499 275807 229527 275835
rect 229561 275807 229589 275835
rect 229623 275807 229651 275835
rect 229437 275745 229465 275773
rect 229499 275745 229527 275773
rect 229561 275745 229589 275773
rect 229623 275745 229651 275773
rect 229437 266931 229465 266959
rect 229499 266931 229527 266959
rect 229561 266931 229589 266959
rect 229623 266931 229651 266959
rect 229437 266869 229465 266897
rect 229499 266869 229527 266897
rect 229561 266869 229589 266897
rect 229623 266869 229651 266897
rect 229437 266807 229465 266835
rect 229499 266807 229527 266835
rect 229561 266807 229589 266835
rect 229623 266807 229651 266835
rect 229437 266745 229465 266773
rect 229499 266745 229527 266773
rect 229561 266745 229589 266773
rect 229623 266745 229651 266773
rect 229437 257931 229465 257959
rect 229499 257931 229527 257959
rect 229561 257931 229589 257959
rect 229623 257931 229651 257959
rect 229437 257869 229465 257897
rect 229499 257869 229527 257897
rect 229561 257869 229589 257897
rect 229623 257869 229651 257897
rect 229437 257807 229465 257835
rect 229499 257807 229527 257835
rect 229561 257807 229589 257835
rect 229623 257807 229651 257835
rect 229437 257745 229465 257773
rect 229499 257745 229527 257773
rect 229561 257745 229589 257773
rect 229623 257745 229651 257773
rect 236577 299162 236605 299190
rect 236639 299162 236667 299190
rect 236701 299162 236729 299190
rect 236763 299162 236791 299190
rect 236577 299100 236605 299128
rect 236639 299100 236667 299128
rect 236701 299100 236729 299128
rect 236763 299100 236791 299128
rect 236577 299038 236605 299066
rect 236639 299038 236667 299066
rect 236701 299038 236729 299066
rect 236763 299038 236791 299066
rect 236577 298976 236605 299004
rect 236639 298976 236667 299004
rect 236701 298976 236729 299004
rect 236763 298976 236791 299004
rect 236577 290931 236605 290959
rect 236639 290931 236667 290959
rect 236701 290931 236729 290959
rect 236763 290931 236791 290959
rect 236577 290869 236605 290897
rect 236639 290869 236667 290897
rect 236701 290869 236729 290897
rect 236763 290869 236791 290897
rect 236577 290807 236605 290835
rect 236639 290807 236667 290835
rect 236701 290807 236729 290835
rect 236763 290807 236791 290835
rect 236577 290745 236605 290773
rect 236639 290745 236667 290773
rect 236701 290745 236729 290773
rect 236763 290745 236791 290773
rect 236577 281931 236605 281959
rect 236639 281931 236667 281959
rect 236701 281931 236729 281959
rect 236763 281931 236791 281959
rect 236577 281869 236605 281897
rect 236639 281869 236667 281897
rect 236701 281869 236729 281897
rect 236763 281869 236791 281897
rect 236577 281807 236605 281835
rect 236639 281807 236667 281835
rect 236701 281807 236729 281835
rect 236763 281807 236791 281835
rect 236577 281745 236605 281773
rect 236639 281745 236667 281773
rect 236701 281745 236729 281773
rect 236763 281745 236791 281773
rect 236577 272931 236605 272959
rect 236639 272931 236667 272959
rect 236701 272931 236729 272959
rect 236763 272931 236791 272959
rect 236577 272869 236605 272897
rect 236639 272869 236667 272897
rect 236701 272869 236729 272897
rect 236763 272869 236791 272897
rect 236577 272807 236605 272835
rect 236639 272807 236667 272835
rect 236701 272807 236729 272835
rect 236763 272807 236791 272835
rect 236577 272745 236605 272773
rect 236639 272745 236667 272773
rect 236701 272745 236729 272773
rect 236763 272745 236791 272773
rect 236577 263931 236605 263959
rect 236639 263931 236667 263959
rect 236701 263931 236729 263959
rect 236763 263931 236791 263959
rect 236577 263869 236605 263897
rect 236639 263869 236667 263897
rect 236701 263869 236729 263897
rect 236763 263869 236791 263897
rect 236577 263807 236605 263835
rect 236639 263807 236667 263835
rect 236701 263807 236729 263835
rect 236763 263807 236791 263835
rect 236577 263745 236605 263773
rect 236639 263745 236667 263773
rect 236701 263745 236729 263773
rect 236763 263745 236791 263773
rect 236577 254931 236605 254959
rect 236639 254931 236667 254959
rect 236701 254931 236729 254959
rect 236763 254931 236791 254959
rect 236577 254869 236605 254897
rect 236639 254869 236667 254897
rect 236701 254869 236729 254897
rect 236763 254869 236791 254897
rect 236577 254807 236605 254835
rect 236639 254807 236667 254835
rect 236701 254807 236729 254835
rect 236763 254807 236791 254835
rect 236577 254745 236605 254773
rect 236639 254745 236667 254773
rect 236701 254745 236729 254773
rect 236763 254745 236791 254773
rect 238437 299642 238465 299670
rect 238499 299642 238527 299670
rect 238561 299642 238589 299670
rect 238623 299642 238651 299670
rect 238437 299580 238465 299608
rect 238499 299580 238527 299608
rect 238561 299580 238589 299608
rect 238623 299580 238651 299608
rect 238437 299518 238465 299546
rect 238499 299518 238527 299546
rect 238561 299518 238589 299546
rect 238623 299518 238651 299546
rect 238437 299456 238465 299484
rect 238499 299456 238527 299484
rect 238561 299456 238589 299484
rect 238623 299456 238651 299484
rect 238437 293931 238465 293959
rect 238499 293931 238527 293959
rect 238561 293931 238589 293959
rect 238623 293931 238651 293959
rect 238437 293869 238465 293897
rect 238499 293869 238527 293897
rect 238561 293869 238589 293897
rect 238623 293869 238651 293897
rect 238437 293807 238465 293835
rect 238499 293807 238527 293835
rect 238561 293807 238589 293835
rect 238623 293807 238651 293835
rect 238437 293745 238465 293773
rect 238499 293745 238527 293773
rect 238561 293745 238589 293773
rect 238623 293745 238651 293773
rect 238437 284931 238465 284959
rect 238499 284931 238527 284959
rect 238561 284931 238589 284959
rect 238623 284931 238651 284959
rect 238437 284869 238465 284897
rect 238499 284869 238527 284897
rect 238561 284869 238589 284897
rect 238623 284869 238651 284897
rect 238437 284807 238465 284835
rect 238499 284807 238527 284835
rect 238561 284807 238589 284835
rect 238623 284807 238651 284835
rect 238437 284745 238465 284773
rect 238499 284745 238527 284773
rect 238561 284745 238589 284773
rect 238623 284745 238651 284773
rect 238437 275931 238465 275959
rect 238499 275931 238527 275959
rect 238561 275931 238589 275959
rect 238623 275931 238651 275959
rect 238437 275869 238465 275897
rect 238499 275869 238527 275897
rect 238561 275869 238589 275897
rect 238623 275869 238651 275897
rect 238437 275807 238465 275835
rect 238499 275807 238527 275835
rect 238561 275807 238589 275835
rect 238623 275807 238651 275835
rect 238437 275745 238465 275773
rect 238499 275745 238527 275773
rect 238561 275745 238589 275773
rect 238623 275745 238651 275773
rect 238437 266931 238465 266959
rect 238499 266931 238527 266959
rect 238561 266931 238589 266959
rect 238623 266931 238651 266959
rect 238437 266869 238465 266897
rect 238499 266869 238527 266897
rect 238561 266869 238589 266897
rect 238623 266869 238651 266897
rect 238437 266807 238465 266835
rect 238499 266807 238527 266835
rect 238561 266807 238589 266835
rect 238623 266807 238651 266835
rect 238437 266745 238465 266773
rect 238499 266745 238527 266773
rect 238561 266745 238589 266773
rect 238623 266745 238651 266773
rect 238437 257931 238465 257959
rect 238499 257931 238527 257959
rect 238561 257931 238589 257959
rect 238623 257931 238651 257959
rect 238437 257869 238465 257897
rect 238499 257869 238527 257897
rect 238561 257869 238589 257897
rect 238623 257869 238651 257897
rect 238437 257807 238465 257835
rect 238499 257807 238527 257835
rect 238561 257807 238589 257835
rect 238623 257807 238651 257835
rect 238437 257745 238465 257773
rect 238499 257745 238527 257773
rect 238561 257745 238589 257773
rect 238623 257745 238651 257773
rect 245577 299162 245605 299190
rect 245639 299162 245667 299190
rect 245701 299162 245729 299190
rect 245763 299162 245791 299190
rect 245577 299100 245605 299128
rect 245639 299100 245667 299128
rect 245701 299100 245729 299128
rect 245763 299100 245791 299128
rect 245577 299038 245605 299066
rect 245639 299038 245667 299066
rect 245701 299038 245729 299066
rect 245763 299038 245791 299066
rect 245577 298976 245605 299004
rect 245639 298976 245667 299004
rect 245701 298976 245729 299004
rect 245763 298976 245791 299004
rect 245577 290931 245605 290959
rect 245639 290931 245667 290959
rect 245701 290931 245729 290959
rect 245763 290931 245791 290959
rect 245577 290869 245605 290897
rect 245639 290869 245667 290897
rect 245701 290869 245729 290897
rect 245763 290869 245791 290897
rect 245577 290807 245605 290835
rect 245639 290807 245667 290835
rect 245701 290807 245729 290835
rect 245763 290807 245791 290835
rect 245577 290745 245605 290773
rect 245639 290745 245667 290773
rect 245701 290745 245729 290773
rect 245763 290745 245791 290773
rect 245577 281931 245605 281959
rect 245639 281931 245667 281959
rect 245701 281931 245729 281959
rect 245763 281931 245791 281959
rect 245577 281869 245605 281897
rect 245639 281869 245667 281897
rect 245701 281869 245729 281897
rect 245763 281869 245791 281897
rect 245577 281807 245605 281835
rect 245639 281807 245667 281835
rect 245701 281807 245729 281835
rect 245763 281807 245791 281835
rect 245577 281745 245605 281773
rect 245639 281745 245667 281773
rect 245701 281745 245729 281773
rect 245763 281745 245791 281773
rect 245577 272931 245605 272959
rect 245639 272931 245667 272959
rect 245701 272931 245729 272959
rect 245763 272931 245791 272959
rect 245577 272869 245605 272897
rect 245639 272869 245667 272897
rect 245701 272869 245729 272897
rect 245763 272869 245791 272897
rect 245577 272807 245605 272835
rect 245639 272807 245667 272835
rect 245701 272807 245729 272835
rect 245763 272807 245791 272835
rect 245577 272745 245605 272773
rect 245639 272745 245667 272773
rect 245701 272745 245729 272773
rect 245763 272745 245791 272773
rect 245577 263931 245605 263959
rect 245639 263931 245667 263959
rect 245701 263931 245729 263959
rect 245763 263931 245791 263959
rect 245577 263869 245605 263897
rect 245639 263869 245667 263897
rect 245701 263869 245729 263897
rect 245763 263869 245791 263897
rect 245577 263807 245605 263835
rect 245639 263807 245667 263835
rect 245701 263807 245729 263835
rect 245763 263807 245791 263835
rect 245577 263745 245605 263773
rect 245639 263745 245667 263773
rect 245701 263745 245729 263773
rect 245763 263745 245791 263773
rect 245577 254931 245605 254959
rect 245639 254931 245667 254959
rect 245701 254931 245729 254959
rect 245763 254931 245791 254959
rect 245577 254869 245605 254897
rect 245639 254869 245667 254897
rect 245701 254869 245729 254897
rect 245763 254869 245791 254897
rect 245577 254807 245605 254835
rect 245639 254807 245667 254835
rect 245701 254807 245729 254835
rect 245763 254807 245791 254835
rect 245577 254745 245605 254773
rect 245639 254745 245667 254773
rect 245701 254745 245729 254773
rect 245763 254745 245791 254773
rect 247437 299642 247465 299670
rect 247499 299642 247527 299670
rect 247561 299642 247589 299670
rect 247623 299642 247651 299670
rect 247437 299580 247465 299608
rect 247499 299580 247527 299608
rect 247561 299580 247589 299608
rect 247623 299580 247651 299608
rect 247437 299518 247465 299546
rect 247499 299518 247527 299546
rect 247561 299518 247589 299546
rect 247623 299518 247651 299546
rect 247437 299456 247465 299484
rect 247499 299456 247527 299484
rect 247561 299456 247589 299484
rect 247623 299456 247651 299484
rect 247437 293931 247465 293959
rect 247499 293931 247527 293959
rect 247561 293931 247589 293959
rect 247623 293931 247651 293959
rect 247437 293869 247465 293897
rect 247499 293869 247527 293897
rect 247561 293869 247589 293897
rect 247623 293869 247651 293897
rect 247437 293807 247465 293835
rect 247499 293807 247527 293835
rect 247561 293807 247589 293835
rect 247623 293807 247651 293835
rect 247437 293745 247465 293773
rect 247499 293745 247527 293773
rect 247561 293745 247589 293773
rect 247623 293745 247651 293773
rect 247437 284931 247465 284959
rect 247499 284931 247527 284959
rect 247561 284931 247589 284959
rect 247623 284931 247651 284959
rect 247437 284869 247465 284897
rect 247499 284869 247527 284897
rect 247561 284869 247589 284897
rect 247623 284869 247651 284897
rect 247437 284807 247465 284835
rect 247499 284807 247527 284835
rect 247561 284807 247589 284835
rect 247623 284807 247651 284835
rect 247437 284745 247465 284773
rect 247499 284745 247527 284773
rect 247561 284745 247589 284773
rect 247623 284745 247651 284773
rect 247437 275931 247465 275959
rect 247499 275931 247527 275959
rect 247561 275931 247589 275959
rect 247623 275931 247651 275959
rect 247437 275869 247465 275897
rect 247499 275869 247527 275897
rect 247561 275869 247589 275897
rect 247623 275869 247651 275897
rect 247437 275807 247465 275835
rect 247499 275807 247527 275835
rect 247561 275807 247589 275835
rect 247623 275807 247651 275835
rect 247437 275745 247465 275773
rect 247499 275745 247527 275773
rect 247561 275745 247589 275773
rect 247623 275745 247651 275773
rect 247437 266931 247465 266959
rect 247499 266931 247527 266959
rect 247561 266931 247589 266959
rect 247623 266931 247651 266959
rect 247437 266869 247465 266897
rect 247499 266869 247527 266897
rect 247561 266869 247589 266897
rect 247623 266869 247651 266897
rect 247437 266807 247465 266835
rect 247499 266807 247527 266835
rect 247561 266807 247589 266835
rect 247623 266807 247651 266835
rect 247437 266745 247465 266773
rect 247499 266745 247527 266773
rect 247561 266745 247589 266773
rect 247623 266745 247651 266773
rect 247437 257931 247465 257959
rect 247499 257931 247527 257959
rect 247561 257931 247589 257959
rect 247623 257931 247651 257959
rect 247437 257869 247465 257897
rect 247499 257869 247527 257897
rect 247561 257869 247589 257897
rect 247623 257869 247651 257897
rect 247437 257807 247465 257835
rect 247499 257807 247527 257835
rect 247561 257807 247589 257835
rect 247623 257807 247651 257835
rect 247437 257745 247465 257773
rect 247499 257745 247527 257773
rect 247561 257745 247589 257773
rect 247623 257745 247651 257773
rect 254577 299162 254605 299190
rect 254639 299162 254667 299190
rect 254701 299162 254729 299190
rect 254763 299162 254791 299190
rect 254577 299100 254605 299128
rect 254639 299100 254667 299128
rect 254701 299100 254729 299128
rect 254763 299100 254791 299128
rect 254577 299038 254605 299066
rect 254639 299038 254667 299066
rect 254701 299038 254729 299066
rect 254763 299038 254791 299066
rect 254577 298976 254605 299004
rect 254639 298976 254667 299004
rect 254701 298976 254729 299004
rect 254763 298976 254791 299004
rect 254577 290931 254605 290959
rect 254639 290931 254667 290959
rect 254701 290931 254729 290959
rect 254763 290931 254791 290959
rect 254577 290869 254605 290897
rect 254639 290869 254667 290897
rect 254701 290869 254729 290897
rect 254763 290869 254791 290897
rect 254577 290807 254605 290835
rect 254639 290807 254667 290835
rect 254701 290807 254729 290835
rect 254763 290807 254791 290835
rect 254577 290745 254605 290773
rect 254639 290745 254667 290773
rect 254701 290745 254729 290773
rect 254763 290745 254791 290773
rect 254577 281931 254605 281959
rect 254639 281931 254667 281959
rect 254701 281931 254729 281959
rect 254763 281931 254791 281959
rect 254577 281869 254605 281897
rect 254639 281869 254667 281897
rect 254701 281869 254729 281897
rect 254763 281869 254791 281897
rect 254577 281807 254605 281835
rect 254639 281807 254667 281835
rect 254701 281807 254729 281835
rect 254763 281807 254791 281835
rect 254577 281745 254605 281773
rect 254639 281745 254667 281773
rect 254701 281745 254729 281773
rect 254763 281745 254791 281773
rect 254577 272931 254605 272959
rect 254639 272931 254667 272959
rect 254701 272931 254729 272959
rect 254763 272931 254791 272959
rect 254577 272869 254605 272897
rect 254639 272869 254667 272897
rect 254701 272869 254729 272897
rect 254763 272869 254791 272897
rect 254577 272807 254605 272835
rect 254639 272807 254667 272835
rect 254701 272807 254729 272835
rect 254763 272807 254791 272835
rect 254577 272745 254605 272773
rect 254639 272745 254667 272773
rect 254701 272745 254729 272773
rect 254763 272745 254791 272773
rect 254577 263931 254605 263959
rect 254639 263931 254667 263959
rect 254701 263931 254729 263959
rect 254763 263931 254791 263959
rect 254577 263869 254605 263897
rect 254639 263869 254667 263897
rect 254701 263869 254729 263897
rect 254763 263869 254791 263897
rect 254577 263807 254605 263835
rect 254639 263807 254667 263835
rect 254701 263807 254729 263835
rect 254763 263807 254791 263835
rect 254577 263745 254605 263773
rect 254639 263745 254667 263773
rect 254701 263745 254729 263773
rect 254763 263745 254791 263773
rect 256437 299642 256465 299670
rect 256499 299642 256527 299670
rect 256561 299642 256589 299670
rect 256623 299642 256651 299670
rect 256437 299580 256465 299608
rect 256499 299580 256527 299608
rect 256561 299580 256589 299608
rect 256623 299580 256651 299608
rect 256437 299518 256465 299546
rect 256499 299518 256527 299546
rect 256561 299518 256589 299546
rect 256623 299518 256651 299546
rect 256437 299456 256465 299484
rect 256499 299456 256527 299484
rect 256561 299456 256589 299484
rect 256623 299456 256651 299484
rect 256437 293931 256465 293959
rect 256499 293931 256527 293959
rect 256561 293931 256589 293959
rect 256623 293931 256651 293959
rect 256437 293869 256465 293897
rect 256499 293869 256527 293897
rect 256561 293869 256589 293897
rect 256623 293869 256651 293897
rect 256437 293807 256465 293835
rect 256499 293807 256527 293835
rect 256561 293807 256589 293835
rect 256623 293807 256651 293835
rect 256437 293745 256465 293773
rect 256499 293745 256527 293773
rect 256561 293745 256589 293773
rect 256623 293745 256651 293773
rect 256437 284931 256465 284959
rect 256499 284931 256527 284959
rect 256561 284931 256589 284959
rect 256623 284931 256651 284959
rect 256437 284869 256465 284897
rect 256499 284869 256527 284897
rect 256561 284869 256589 284897
rect 256623 284869 256651 284897
rect 256437 284807 256465 284835
rect 256499 284807 256527 284835
rect 256561 284807 256589 284835
rect 256623 284807 256651 284835
rect 256437 284745 256465 284773
rect 256499 284745 256527 284773
rect 256561 284745 256589 284773
rect 256623 284745 256651 284773
rect 256437 275931 256465 275959
rect 256499 275931 256527 275959
rect 256561 275931 256589 275959
rect 256623 275931 256651 275959
rect 256437 275869 256465 275897
rect 256499 275869 256527 275897
rect 256561 275869 256589 275897
rect 256623 275869 256651 275897
rect 256437 275807 256465 275835
rect 256499 275807 256527 275835
rect 256561 275807 256589 275835
rect 256623 275807 256651 275835
rect 256437 275745 256465 275773
rect 256499 275745 256527 275773
rect 256561 275745 256589 275773
rect 256623 275745 256651 275773
rect 256437 266931 256465 266959
rect 256499 266931 256527 266959
rect 256561 266931 256589 266959
rect 256623 266931 256651 266959
rect 256437 266869 256465 266897
rect 256499 266869 256527 266897
rect 256561 266869 256589 266897
rect 256623 266869 256651 266897
rect 256437 266807 256465 266835
rect 256499 266807 256527 266835
rect 256561 266807 256589 266835
rect 256623 266807 256651 266835
rect 256437 266745 256465 266773
rect 256499 266745 256527 266773
rect 256561 266745 256589 266773
rect 256623 266745 256651 266773
rect 256437 257931 256465 257959
rect 256499 257931 256527 257959
rect 256561 257931 256589 257959
rect 256623 257931 256651 257959
rect 256437 257869 256465 257897
rect 256499 257869 256527 257897
rect 256561 257869 256589 257897
rect 256623 257869 256651 257897
rect 256437 257807 256465 257835
rect 256499 257807 256527 257835
rect 256561 257807 256589 257835
rect 256623 257807 256651 257835
rect 256437 257745 256465 257773
rect 256499 257745 256527 257773
rect 256561 257745 256589 257773
rect 256623 257745 256651 257773
rect 254577 254931 254605 254959
rect 254639 254931 254667 254959
rect 254701 254931 254729 254959
rect 254763 254931 254791 254959
rect 254577 254869 254605 254897
rect 254639 254869 254667 254897
rect 254701 254869 254729 254897
rect 254763 254869 254791 254897
rect 254577 254807 254605 254835
rect 254639 254807 254667 254835
rect 254701 254807 254729 254835
rect 254763 254807 254791 254835
rect 254577 254745 254605 254773
rect 254639 254745 254667 254773
rect 254701 254745 254729 254773
rect 254763 254745 254791 254773
rect 31437 248931 31465 248959
rect 31499 248931 31527 248959
rect 31561 248931 31589 248959
rect 31623 248931 31651 248959
rect 31437 248869 31465 248897
rect 31499 248869 31527 248897
rect 31561 248869 31589 248897
rect 31623 248869 31651 248897
rect 31437 248807 31465 248835
rect 31499 248807 31527 248835
rect 31561 248807 31589 248835
rect 31623 248807 31651 248835
rect 31437 248745 31465 248773
rect 31499 248745 31527 248773
rect 31561 248745 31589 248773
rect 31623 248745 31651 248773
rect 40299 248931 40327 248959
rect 40361 248931 40389 248959
rect 40299 248869 40327 248897
rect 40361 248869 40389 248897
rect 40299 248807 40327 248835
rect 40361 248807 40389 248835
rect 40299 248745 40327 248773
rect 40361 248745 40389 248773
rect 55659 248931 55687 248959
rect 55721 248931 55749 248959
rect 55659 248869 55687 248897
rect 55721 248869 55749 248897
rect 55659 248807 55687 248835
rect 55721 248807 55749 248835
rect 55659 248745 55687 248773
rect 55721 248745 55749 248773
rect 71019 248931 71047 248959
rect 71081 248931 71109 248959
rect 71019 248869 71047 248897
rect 71081 248869 71109 248897
rect 71019 248807 71047 248835
rect 71081 248807 71109 248835
rect 71019 248745 71047 248773
rect 71081 248745 71109 248773
rect 86379 248931 86407 248959
rect 86441 248931 86469 248959
rect 86379 248869 86407 248897
rect 86441 248869 86469 248897
rect 86379 248807 86407 248835
rect 86441 248807 86469 248835
rect 86379 248745 86407 248773
rect 86441 248745 86469 248773
rect 101739 248931 101767 248959
rect 101801 248931 101829 248959
rect 101739 248869 101767 248897
rect 101801 248869 101829 248897
rect 101739 248807 101767 248835
rect 101801 248807 101829 248835
rect 101739 248745 101767 248773
rect 101801 248745 101829 248773
rect 117099 248931 117127 248959
rect 117161 248931 117189 248959
rect 117099 248869 117127 248897
rect 117161 248869 117189 248897
rect 117099 248807 117127 248835
rect 117161 248807 117189 248835
rect 117099 248745 117127 248773
rect 117161 248745 117189 248773
rect 132459 248931 132487 248959
rect 132521 248931 132549 248959
rect 132459 248869 132487 248897
rect 132521 248869 132549 248897
rect 132459 248807 132487 248835
rect 132521 248807 132549 248835
rect 132459 248745 132487 248773
rect 132521 248745 132549 248773
rect 147819 248931 147847 248959
rect 147881 248931 147909 248959
rect 147819 248869 147847 248897
rect 147881 248869 147909 248897
rect 147819 248807 147847 248835
rect 147881 248807 147909 248835
rect 147819 248745 147847 248773
rect 147881 248745 147909 248773
rect 163179 248931 163207 248959
rect 163241 248931 163269 248959
rect 163179 248869 163207 248897
rect 163241 248869 163269 248897
rect 163179 248807 163207 248835
rect 163241 248807 163269 248835
rect 163179 248745 163207 248773
rect 163241 248745 163269 248773
rect 178539 248931 178567 248959
rect 178601 248931 178629 248959
rect 178539 248869 178567 248897
rect 178601 248869 178629 248897
rect 178539 248807 178567 248835
rect 178601 248807 178629 248835
rect 178539 248745 178567 248773
rect 178601 248745 178629 248773
rect 193899 248931 193927 248959
rect 193961 248931 193989 248959
rect 193899 248869 193927 248897
rect 193961 248869 193989 248897
rect 193899 248807 193927 248835
rect 193961 248807 193989 248835
rect 193899 248745 193927 248773
rect 193961 248745 193989 248773
rect 209259 248931 209287 248959
rect 209321 248931 209349 248959
rect 209259 248869 209287 248897
rect 209321 248869 209349 248897
rect 209259 248807 209287 248835
rect 209321 248807 209349 248835
rect 209259 248745 209287 248773
rect 209321 248745 209349 248773
rect 224619 248931 224647 248959
rect 224681 248931 224709 248959
rect 224619 248869 224647 248897
rect 224681 248869 224709 248897
rect 224619 248807 224647 248835
rect 224681 248807 224709 248835
rect 224619 248745 224647 248773
rect 224681 248745 224709 248773
rect 239979 248931 240007 248959
rect 240041 248931 240069 248959
rect 239979 248869 240007 248897
rect 240041 248869 240069 248897
rect 239979 248807 240007 248835
rect 240041 248807 240069 248835
rect 239979 248745 240007 248773
rect 240041 248745 240069 248773
rect 32619 245931 32647 245959
rect 32681 245931 32709 245959
rect 32619 245869 32647 245897
rect 32681 245869 32709 245897
rect 32619 245807 32647 245835
rect 32681 245807 32709 245835
rect 32619 245745 32647 245773
rect 32681 245745 32709 245773
rect 47979 245931 48007 245959
rect 48041 245931 48069 245959
rect 47979 245869 48007 245897
rect 48041 245869 48069 245897
rect 47979 245807 48007 245835
rect 48041 245807 48069 245835
rect 47979 245745 48007 245773
rect 48041 245745 48069 245773
rect 63339 245931 63367 245959
rect 63401 245931 63429 245959
rect 63339 245869 63367 245897
rect 63401 245869 63429 245897
rect 63339 245807 63367 245835
rect 63401 245807 63429 245835
rect 63339 245745 63367 245773
rect 63401 245745 63429 245773
rect 78699 245931 78727 245959
rect 78761 245931 78789 245959
rect 78699 245869 78727 245897
rect 78761 245869 78789 245897
rect 78699 245807 78727 245835
rect 78761 245807 78789 245835
rect 78699 245745 78727 245773
rect 78761 245745 78789 245773
rect 94059 245931 94087 245959
rect 94121 245931 94149 245959
rect 94059 245869 94087 245897
rect 94121 245869 94149 245897
rect 94059 245807 94087 245835
rect 94121 245807 94149 245835
rect 94059 245745 94087 245773
rect 94121 245745 94149 245773
rect 109419 245931 109447 245959
rect 109481 245931 109509 245959
rect 109419 245869 109447 245897
rect 109481 245869 109509 245897
rect 109419 245807 109447 245835
rect 109481 245807 109509 245835
rect 109419 245745 109447 245773
rect 109481 245745 109509 245773
rect 124779 245931 124807 245959
rect 124841 245931 124869 245959
rect 124779 245869 124807 245897
rect 124841 245869 124869 245897
rect 124779 245807 124807 245835
rect 124841 245807 124869 245835
rect 124779 245745 124807 245773
rect 124841 245745 124869 245773
rect 140139 245931 140167 245959
rect 140201 245931 140229 245959
rect 140139 245869 140167 245897
rect 140201 245869 140229 245897
rect 140139 245807 140167 245835
rect 140201 245807 140229 245835
rect 140139 245745 140167 245773
rect 140201 245745 140229 245773
rect 155499 245931 155527 245959
rect 155561 245931 155589 245959
rect 155499 245869 155527 245897
rect 155561 245869 155589 245897
rect 155499 245807 155527 245835
rect 155561 245807 155589 245835
rect 155499 245745 155527 245773
rect 155561 245745 155589 245773
rect 170859 245931 170887 245959
rect 170921 245931 170949 245959
rect 170859 245869 170887 245897
rect 170921 245869 170949 245897
rect 170859 245807 170887 245835
rect 170921 245807 170949 245835
rect 170859 245745 170887 245773
rect 170921 245745 170949 245773
rect 186219 245931 186247 245959
rect 186281 245931 186309 245959
rect 186219 245869 186247 245897
rect 186281 245869 186309 245897
rect 186219 245807 186247 245835
rect 186281 245807 186309 245835
rect 186219 245745 186247 245773
rect 186281 245745 186309 245773
rect 201579 245931 201607 245959
rect 201641 245931 201669 245959
rect 201579 245869 201607 245897
rect 201641 245869 201669 245897
rect 201579 245807 201607 245835
rect 201641 245807 201669 245835
rect 201579 245745 201607 245773
rect 201641 245745 201669 245773
rect 216939 245931 216967 245959
rect 217001 245931 217029 245959
rect 216939 245869 216967 245897
rect 217001 245869 217029 245897
rect 216939 245807 216967 245835
rect 217001 245807 217029 245835
rect 216939 245745 216967 245773
rect 217001 245745 217029 245773
rect 232299 245931 232327 245959
rect 232361 245931 232389 245959
rect 232299 245869 232327 245897
rect 232361 245869 232389 245897
rect 232299 245807 232327 245835
rect 232361 245807 232389 245835
rect 232299 245745 232327 245773
rect 232361 245745 232389 245773
rect 247659 245931 247687 245959
rect 247721 245931 247749 245959
rect 247659 245869 247687 245897
rect 247721 245869 247749 245897
rect 247659 245807 247687 245835
rect 247721 245807 247749 245835
rect 247659 245745 247687 245773
rect 247721 245745 247749 245773
rect 254577 245931 254605 245959
rect 254639 245931 254667 245959
rect 254701 245931 254729 245959
rect 254763 245931 254791 245959
rect 254577 245869 254605 245897
rect 254639 245869 254667 245897
rect 254701 245869 254729 245897
rect 254763 245869 254791 245897
rect 254577 245807 254605 245835
rect 254639 245807 254667 245835
rect 254701 245807 254729 245835
rect 254763 245807 254791 245835
rect 254577 245745 254605 245773
rect 254639 245745 254667 245773
rect 254701 245745 254729 245773
rect 254763 245745 254791 245773
rect 31437 239931 31465 239959
rect 31499 239931 31527 239959
rect 31561 239931 31589 239959
rect 31623 239931 31651 239959
rect 31437 239869 31465 239897
rect 31499 239869 31527 239897
rect 31561 239869 31589 239897
rect 31623 239869 31651 239897
rect 31437 239807 31465 239835
rect 31499 239807 31527 239835
rect 31561 239807 31589 239835
rect 31623 239807 31651 239835
rect 31437 239745 31465 239773
rect 31499 239745 31527 239773
rect 31561 239745 31589 239773
rect 31623 239745 31651 239773
rect 40299 239931 40327 239959
rect 40361 239931 40389 239959
rect 40299 239869 40327 239897
rect 40361 239869 40389 239897
rect 40299 239807 40327 239835
rect 40361 239807 40389 239835
rect 40299 239745 40327 239773
rect 40361 239745 40389 239773
rect 55659 239931 55687 239959
rect 55721 239931 55749 239959
rect 55659 239869 55687 239897
rect 55721 239869 55749 239897
rect 55659 239807 55687 239835
rect 55721 239807 55749 239835
rect 55659 239745 55687 239773
rect 55721 239745 55749 239773
rect 71019 239931 71047 239959
rect 71081 239931 71109 239959
rect 71019 239869 71047 239897
rect 71081 239869 71109 239897
rect 71019 239807 71047 239835
rect 71081 239807 71109 239835
rect 71019 239745 71047 239773
rect 71081 239745 71109 239773
rect 86379 239931 86407 239959
rect 86441 239931 86469 239959
rect 86379 239869 86407 239897
rect 86441 239869 86469 239897
rect 86379 239807 86407 239835
rect 86441 239807 86469 239835
rect 86379 239745 86407 239773
rect 86441 239745 86469 239773
rect 101739 239931 101767 239959
rect 101801 239931 101829 239959
rect 101739 239869 101767 239897
rect 101801 239869 101829 239897
rect 101739 239807 101767 239835
rect 101801 239807 101829 239835
rect 101739 239745 101767 239773
rect 101801 239745 101829 239773
rect 117099 239931 117127 239959
rect 117161 239931 117189 239959
rect 117099 239869 117127 239897
rect 117161 239869 117189 239897
rect 117099 239807 117127 239835
rect 117161 239807 117189 239835
rect 117099 239745 117127 239773
rect 117161 239745 117189 239773
rect 132459 239931 132487 239959
rect 132521 239931 132549 239959
rect 132459 239869 132487 239897
rect 132521 239869 132549 239897
rect 132459 239807 132487 239835
rect 132521 239807 132549 239835
rect 132459 239745 132487 239773
rect 132521 239745 132549 239773
rect 147819 239931 147847 239959
rect 147881 239931 147909 239959
rect 147819 239869 147847 239897
rect 147881 239869 147909 239897
rect 147819 239807 147847 239835
rect 147881 239807 147909 239835
rect 147819 239745 147847 239773
rect 147881 239745 147909 239773
rect 163179 239931 163207 239959
rect 163241 239931 163269 239959
rect 163179 239869 163207 239897
rect 163241 239869 163269 239897
rect 163179 239807 163207 239835
rect 163241 239807 163269 239835
rect 163179 239745 163207 239773
rect 163241 239745 163269 239773
rect 178539 239931 178567 239959
rect 178601 239931 178629 239959
rect 178539 239869 178567 239897
rect 178601 239869 178629 239897
rect 178539 239807 178567 239835
rect 178601 239807 178629 239835
rect 178539 239745 178567 239773
rect 178601 239745 178629 239773
rect 193899 239931 193927 239959
rect 193961 239931 193989 239959
rect 193899 239869 193927 239897
rect 193961 239869 193989 239897
rect 193899 239807 193927 239835
rect 193961 239807 193989 239835
rect 193899 239745 193927 239773
rect 193961 239745 193989 239773
rect 209259 239931 209287 239959
rect 209321 239931 209349 239959
rect 209259 239869 209287 239897
rect 209321 239869 209349 239897
rect 209259 239807 209287 239835
rect 209321 239807 209349 239835
rect 209259 239745 209287 239773
rect 209321 239745 209349 239773
rect 224619 239931 224647 239959
rect 224681 239931 224709 239959
rect 224619 239869 224647 239897
rect 224681 239869 224709 239897
rect 224619 239807 224647 239835
rect 224681 239807 224709 239835
rect 224619 239745 224647 239773
rect 224681 239745 224709 239773
rect 239979 239931 240007 239959
rect 240041 239931 240069 239959
rect 239979 239869 240007 239897
rect 240041 239869 240069 239897
rect 239979 239807 240007 239835
rect 240041 239807 240069 239835
rect 239979 239745 240007 239773
rect 240041 239745 240069 239773
rect 32619 236931 32647 236959
rect 32681 236931 32709 236959
rect 32619 236869 32647 236897
rect 32681 236869 32709 236897
rect 32619 236807 32647 236835
rect 32681 236807 32709 236835
rect 32619 236745 32647 236773
rect 32681 236745 32709 236773
rect 47979 236931 48007 236959
rect 48041 236931 48069 236959
rect 47979 236869 48007 236897
rect 48041 236869 48069 236897
rect 47979 236807 48007 236835
rect 48041 236807 48069 236835
rect 47979 236745 48007 236773
rect 48041 236745 48069 236773
rect 63339 236931 63367 236959
rect 63401 236931 63429 236959
rect 63339 236869 63367 236897
rect 63401 236869 63429 236897
rect 63339 236807 63367 236835
rect 63401 236807 63429 236835
rect 63339 236745 63367 236773
rect 63401 236745 63429 236773
rect 78699 236931 78727 236959
rect 78761 236931 78789 236959
rect 78699 236869 78727 236897
rect 78761 236869 78789 236897
rect 78699 236807 78727 236835
rect 78761 236807 78789 236835
rect 78699 236745 78727 236773
rect 78761 236745 78789 236773
rect 94059 236931 94087 236959
rect 94121 236931 94149 236959
rect 94059 236869 94087 236897
rect 94121 236869 94149 236897
rect 94059 236807 94087 236835
rect 94121 236807 94149 236835
rect 94059 236745 94087 236773
rect 94121 236745 94149 236773
rect 109419 236931 109447 236959
rect 109481 236931 109509 236959
rect 109419 236869 109447 236897
rect 109481 236869 109509 236897
rect 109419 236807 109447 236835
rect 109481 236807 109509 236835
rect 109419 236745 109447 236773
rect 109481 236745 109509 236773
rect 124779 236931 124807 236959
rect 124841 236931 124869 236959
rect 124779 236869 124807 236897
rect 124841 236869 124869 236897
rect 124779 236807 124807 236835
rect 124841 236807 124869 236835
rect 124779 236745 124807 236773
rect 124841 236745 124869 236773
rect 140139 236931 140167 236959
rect 140201 236931 140229 236959
rect 140139 236869 140167 236897
rect 140201 236869 140229 236897
rect 140139 236807 140167 236835
rect 140201 236807 140229 236835
rect 140139 236745 140167 236773
rect 140201 236745 140229 236773
rect 155499 236931 155527 236959
rect 155561 236931 155589 236959
rect 155499 236869 155527 236897
rect 155561 236869 155589 236897
rect 155499 236807 155527 236835
rect 155561 236807 155589 236835
rect 155499 236745 155527 236773
rect 155561 236745 155589 236773
rect 170859 236931 170887 236959
rect 170921 236931 170949 236959
rect 170859 236869 170887 236897
rect 170921 236869 170949 236897
rect 170859 236807 170887 236835
rect 170921 236807 170949 236835
rect 170859 236745 170887 236773
rect 170921 236745 170949 236773
rect 186219 236931 186247 236959
rect 186281 236931 186309 236959
rect 186219 236869 186247 236897
rect 186281 236869 186309 236897
rect 186219 236807 186247 236835
rect 186281 236807 186309 236835
rect 186219 236745 186247 236773
rect 186281 236745 186309 236773
rect 201579 236931 201607 236959
rect 201641 236931 201669 236959
rect 201579 236869 201607 236897
rect 201641 236869 201669 236897
rect 201579 236807 201607 236835
rect 201641 236807 201669 236835
rect 201579 236745 201607 236773
rect 201641 236745 201669 236773
rect 216939 236931 216967 236959
rect 217001 236931 217029 236959
rect 216939 236869 216967 236897
rect 217001 236869 217029 236897
rect 216939 236807 216967 236835
rect 217001 236807 217029 236835
rect 216939 236745 216967 236773
rect 217001 236745 217029 236773
rect 232299 236931 232327 236959
rect 232361 236931 232389 236959
rect 232299 236869 232327 236897
rect 232361 236869 232389 236897
rect 232299 236807 232327 236835
rect 232361 236807 232389 236835
rect 232299 236745 232327 236773
rect 232361 236745 232389 236773
rect 247659 236931 247687 236959
rect 247721 236931 247749 236959
rect 247659 236869 247687 236897
rect 247721 236869 247749 236897
rect 247659 236807 247687 236835
rect 247721 236807 247749 236835
rect 247659 236745 247687 236773
rect 247721 236745 247749 236773
rect 254577 236931 254605 236959
rect 254639 236931 254667 236959
rect 254701 236931 254729 236959
rect 254763 236931 254791 236959
rect 254577 236869 254605 236897
rect 254639 236869 254667 236897
rect 254701 236869 254729 236897
rect 254763 236869 254791 236897
rect 254577 236807 254605 236835
rect 254639 236807 254667 236835
rect 254701 236807 254729 236835
rect 254763 236807 254791 236835
rect 254577 236745 254605 236773
rect 254639 236745 254667 236773
rect 254701 236745 254729 236773
rect 254763 236745 254791 236773
rect 31437 230931 31465 230959
rect 31499 230931 31527 230959
rect 31561 230931 31589 230959
rect 31623 230931 31651 230959
rect 31437 230869 31465 230897
rect 31499 230869 31527 230897
rect 31561 230869 31589 230897
rect 31623 230869 31651 230897
rect 31437 230807 31465 230835
rect 31499 230807 31527 230835
rect 31561 230807 31589 230835
rect 31623 230807 31651 230835
rect 31437 230745 31465 230773
rect 31499 230745 31527 230773
rect 31561 230745 31589 230773
rect 31623 230745 31651 230773
rect 40299 230931 40327 230959
rect 40361 230931 40389 230959
rect 40299 230869 40327 230897
rect 40361 230869 40389 230897
rect 40299 230807 40327 230835
rect 40361 230807 40389 230835
rect 40299 230745 40327 230773
rect 40361 230745 40389 230773
rect 55659 230931 55687 230959
rect 55721 230931 55749 230959
rect 55659 230869 55687 230897
rect 55721 230869 55749 230897
rect 55659 230807 55687 230835
rect 55721 230807 55749 230835
rect 55659 230745 55687 230773
rect 55721 230745 55749 230773
rect 71019 230931 71047 230959
rect 71081 230931 71109 230959
rect 71019 230869 71047 230897
rect 71081 230869 71109 230897
rect 71019 230807 71047 230835
rect 71081 230807 71109 230835
rect 71019 230745 71047 230773
rect 71081 230745 71109 230773
rect 86379 230931 86407 230959
rect 86441 230931 86469 230959
rect 86379 230869 86407 230897
rect 86441 230869 86469 230897
rect 86379 230807 86407 230835
rect 86441 230807 86469 230835
rect 86379 230745 86407 230773
rect 86441 230745 86469 230773
rect 101739 230931 101767 230959
rect 101801 230931 101829 230959
rect 101739 230869 101767 230897
rect 101801 230869 101829 230897
rect 101739 230807 101767 230835
rect 101801 230807 101829 230835
rect 101739 230745 101767 230773
rect 101801 230745 101829 230773
rect 117099 230931 117127 230959
rect 117161 230931 117189 230959
rect 117099 230869 117127 230897
rect 117161 230869 117189 230897
rect 117099 230807 117127 230835
rect 117161 230807 117189 230835
rect 117099 230745 117127 230773
rect 117161 230745 117189 230773
rect 132459 230931 132487 230959
rect 132521 230931 132549 230959
rect 132459 230869 132487 230897
rect 132521 230869 132549 230897
rect 132459 230807 132487 230835
rect 132521 230807 132549 230835
rect 132459 230745 132487 230773
rect 132521 230745 132549 230773
rect 147819 230931 147847 230959
rect 147881 230931 147909 230959
rect 147819 230869 147847 230897
rect 147881 230869 147909 230897
rect 147819 230807 147847 230835
rect 147881 230807 147909 230835
rect 147819 230745 147847 230773
rect 147881 230745 147909 230773
rect 163179 230931 163207 230959
rect 163241 230931 163269 230959
rect 163179 230869 163207 230897
rect 163241 230869 163269 230897
rect 163179 230807 163207 230835
rect 163241 230807 163269 230835
rect 163179 230745 163207 230773
rect 163241 230745 163269 230773
rect 178539 230931 178567 230959
rect 178601 230931 178629 230959
rect 178539 230869 178567 230897
rect 178601 230869 178629 230897
rect 178539 230807 178567 230835
rect 178601 230807 178629 230835
rect 178539 230745 178567 230773
rect 178601 230745 178629 230773
rect 193899 230931 193927 230959
rect 193961 230931 193989 230959
rect 193899 230869 193927 230897
rect 193961 230869 193989 230897
rect 193899 230807 193927 230835
rect 193961 230807 193989 230835
rect 193899 230745 193927 230773
rect 193961 230745 193989 230773
rect 209259 230931 209287 230959
rect 209321 230931 209349 230959
rect 209259 230869 209287 230897
rect 209321 230869 209349 230897
rect 209259 230807 209287 230835
rect 209321 230807 209349 230835
rect 209259 230745 209287 230773
rect 209321 230745 209349 230773
rect 224619 230931 224647 230959
rect 224681 230931 224709 230959
rect 224619 230869 224647 230897
rect 224681 230869 224709 230897
rect 224619 230807 224647 230835
rect 224681 230807 224709 230835
rect 224619 230745 224647 230773
rect 224681 230745 224709 230773
rect 239979 230931 240007 230959
rect 240041 230931 240069 230959
rect 239979 230869 240007 230897
rect 240041 230869 240069 230897
rect 239979 230807 240007 230835
rect 240041 230807 240069 230835
rect 239979 230745 240007 230773
rect 240041 230745 240069 230773
rect 32619 227931 32647 227959
rect 32681 227931 32709 227959
rect 32619 227869 32647 227897
rect 32681 227869 32709 227897
rect 32619 227807 32647 227835
rect 32681 227807 32709 227835
rect 32619 227745 32647 227773
rect 32681 227745 32709 227773
rect 47979 227931 48007 227959
rect 48041 227931 48069 227959
rect 47979 227869 48007 227897
rect 48041 227869 48069 227897
rect 47979 227807 48007 227835
rect 48041 227807 48069 227835
rect 47979 227745 48007 227773
rect 48041 227745 48069 227773
rect 63339 227931 63367 227959
rect 63401 227931 63429 227959
rect 63339 227869 63367 227897
rect 63401 227869 63429 227897
rect 63339 227807 63367 227835
rect 63401 227807 63429 227835
rect 63339 227745 63367 227773
rect 63401 227745 63429 227773
rect 78699 227931 78727 227959
rect 78761 227931 78789 227959
rect 78699 227869 78727 227897
rect 78761 227869 78789 227897
rect 78699 227807 78727 227835
rect 78761 227807 78789 227835
rect 78699 227745 78727 227773
rect 78761 227745 78789 227773
rect 94059 227931 94087 227959
rect 94121 227931 94149 227959
rect 94059 227869 94087 227897
rect 94121 227869 94149 227897
rect 94059 227807 94087 227835
rect 94121 227807 94149 227835
rect 94059 227745 94087 227773
rect 94121 227745 94149 227773
rect 109419 227931 109447 227959
rect 109481 227931 109509 227959
rect 109419 227869 109447 227897
rect 109481 227869 109509 227897
rect 109419 227807 109447 227835
rect 109481 227807 109509 227835
rect 109419 227745 109447 227773
rect 109481 227745 109509 227773
rect 124779 227931 124807 227959
rect 124841 227931 124869 227959
rect 124779 227869 124807 227897
rect 124841 227869 124869 227897
rect 124779 227807 124807 227835
rect 124841 227807 124869 227835
rect 124779 227745 124807 227773
rect 124841 227745 124869 227773
rect 140139 227931 140167 227959
rect 140201 227931 140229 227959
rect 140139 227869 140167 227897
rect 140201 227869 140229 227897
rect 140139 227807 140167 227835
rect 140201 227807 140229 227835
rect 140139 227745 140167 227773
rect 140201 227745 140229 227773
rect 155499 227931 155527 227959
rect 155561 227931 155589 227959
rect 155499 227869 155527 227897
rect 155561 227869 155589 227897
rect 155499 227807 155527 227835
rect 155561 227807 155589 227835
rect 155499 227745 155527 227773
rect 155561 227745 155589 227773
rect 170859 227931 170887 227959
rect 170921 227931 170949 227959
rect 170859 227869 170887 227897
rect 170921 227869 170949 227897
rect 170859 227807 170887 227835
rect 170921 227807 170949 227835
rect 170859 227745 170887 227773
rect 170921 227745 170949 227773
rect 186219 227931 186247 227959
rect 186281 227931 186309 227959
rect 186219 227869 186247 227897
rect 186281 227869 186309 227897
rect 186219 227807 186247 227835
rect 186281 227807 186309 227835
rect 186219 227745 186247 227773
rect 186281 227745 186309 227773
rect 201579 227931 201607 227959
rect 201641 227931 201669 227959
rect 201579 227869 201607 227897
rect 201641 227869 201669 227897
rect 201579 227807 201607 227835
rect 201641 227807 201669 227835
rect 201579 227745 201607 227773
rect 201641 227745 201669 227773
rect 216939 227931 216967 227959
rect 217001 227931 217029 227959
rect 216939 227869 216967 227897
rect 217001 227869 217029 227897
rect 216939 227807 216967 227835
rect 217001 227807 217029 227835
rect 216939 227745 216967 227773
rect 217001 227745 217029 227773
rect 232299 227931 232327 227959
rect 232361 227931 232389 227959
rect 232299 227869 232327 227897
rect 232361 227869 232389 227897
rect 232299 227807 232327 227835
rect 232361 227807 232389 227835
rect 232299 227745 232327 227773
rect 232361 227745 232389 227773
rect 247659 227931 247687 227959
rect 247721 227931 247749 227959
rect 247659 227869 247687 227897
rect 247721 227869 247749 227897
rect 247659 227807 247687 227835
rect 247721 227807 247749 227835
rect 247659 227745 247687 227773
rect 247721 227745 247749 227773
rect 254577 227931 254605 227959
rect 254639 227931 254667 227959
rect 254701 227931 254729 227959
rect 254763 227931 254791 227959
rect 254577 227869 254605 227897
rect 254639 227869 254667 227897
rect 254701 227869 254729 227897
rect 254763 227869 254791 227897
rect 254577 227807 254605 227835
rect 254639 227807 254667 227835
rect 254701 227807 254729 227835
rect 254763 227807 254791 227835
rect 254577 227745 254605 227773
rect 254639 227745 254667 227773
rect 254701 227745 254729 227773
rect 254763 227745 254791 227773
rect 31437 221931 31465 221959
rect 31499 221931 31527 221959
rect 31561 221931 31589 221959
rect 31623 221931 31651 221959
rect 31437 221869 31465 221897
rect 31499 221869 31527 221897
rect 31561 221869 31589 221897
rect 31623 221869 31651 221897
rect 31437 221807 31465 221835
rect 31499 221807 31527 221835
rect 31561 221807 31589 221835
rect 31623 221807 31651 221835
rect 31437 221745 31465 221773
rect 31499 221745 31527 221773
rect 31561 221745 31589 221773
rect 31623 221745 31651 221773
rect 40299 221931 40327 221959
rect 40361 221931 40389 221959
rect 40299 221869 40327 221897
rect 40361 221869 40389 221897
rect 40299 221807 40327 221835
rect 40361 221807 40389 221835
rect 40299 221745 40327 221773
rect 40361 221745 40389 221773
rect 55659 221931 55687 221959
rect 55721 221931 55749 221959
rect 55659 221869 55687 221897
rect 55721 221869 55749 221897
rect 55659 221807 55687 221835
rect 55721 221807 55749 221835
rect 55659 221745 55687 221773
rect 55721 221745 55749 221773
rect 71019 221931 71047 221959
rect 71081 221931 71109 221959
rect 71019 221869 71047 221897
rect 71081 221869 71109 221897
rect 71019 221807 71047 221835
rect 71081 221807 71109 221835
rect 71019 221745 71047 221773
rect 71081 221745 71109 221773
rect 86379 221931 86407 221959
rect 86441 221931 86469 221959
rect 86379 221869 86407 221897
rect 86441 221869 86469 221897
rect 86379 221807 86407 221835
rect 86441 221807 86469 221835
rect 86379 221745 86407 221773
rect 86441 221745 86469 221773
rect 101739 221931 101767 221959
rect 101801 221931 101829 221959
rect 101739 221869 101767 221897
rect 101801 221869 101829 221897
rect 101739 221807 101767 221835
rect 101801 221807 101829 221835
rect 101739 221745 101767 221773
rect 101801 221745 101829 221773
rect 117099 221931 117127 221959
rect 117161 221931 117189 221959
rect 117099 221869 117127 221897
rect 117161 221869 117189 221897
rect 117099 221807 117127 221835
rect 117161 221807 117189 221835
rect 117099 221745 117127 221773
rect 117161 221745 117189 221773
rect 132459 221931 132487 221959
rect 132521 221931 132549 221959
rect 132459 221869 132487 221897
rect 132521 221869 132549 221897
rect 132459 221807 132487 221835
rect 132521 221807 132549 221835
rect 132459 221745 132487 221773
rect 132521 221745 132549 221773
rect 147819 221931 147847 221959
rect 147881 221931 147909 221959
rect 147819 221869 147847 221897
rect 147881 221869 147909 221897
rect 147819 221807 147847 221835
rect 147881 221807 147909 221835
rect 147819 221745 147847 221773
rect 147881 221745 147909 221773
rect 163179 221931 163207 221959
rect 163241 221931 163269 221959
rect 163179 221869 163207 221897
rect 163241 221869 163269 221897
rect 163179 221807 163207 221835
rect 163241 221807 163269 221835
rect 163179 221745 163207 221773
rect 163241 221745 163269 221773
rect 178539 221931 178567 221959
rect 178601 221931 178629 221959
rect 178539 221869 178567 221897
rect 178601 221869 178629 221897
rect 178539 221807 178567 221835
rect 178601 221807 178629 221835
rect 178539 221745 178567 221773
rect 178601 221745 178629 221773
rect 193899 221931 193927 221959
rect 193961 221931 193989 221959
rect 193899 221869 193927 221897
rect 193961 221869 193989 221897
rect 193899 221807 193927 221835
rect 193961 221807 193989 221835
rect 193899 221745 193927 221773
rect 193961 221745 193989 221773
rect 209259 221931 209287 221959
rect 209321 221931 209349 221959
rect 209259 221869 209287 221897
rect 209321 221869 209349 221897
rect 209259 221807 209287 221835
rect 209321 221807 209349 221835
rect 209259 221745 209287 221773
rect 209321 221745 209349 221773
rect 224619 221931 224647 221959
rect 224681 221931 224709 221959
rect 224619 221869 224647 221897
rect 224681 221869 224709 221897
rect 224619 221807 224647 221835
rect 224681 221807 224709 221835
rect 224619 221745 224647 221773
rect 224681 221745 224709 221773
rect 239979 221931 240007 221959
rect 240041 221931 240069 221959
rect 239979 221869 240007 221897
rect 240041 221869 240069 221897
rect 239979 221807 240007 221835
rect 240041 221807 240069 221835
rect 239979 221745 240007 221773
rect 240041 221745 240069 221773
rect 32619 218931 32647 218959
rect 32681 218931 32709 218959
rect 32619 218869 32647 218897
rect 32681 218869 32709 218897
rect 32619 218807 32647 218835
rect 32681 218807 32709 218835
rect 32619 218745 32647 218773
rect 32681 218745 32709 218773
rect 47979 218931 48007 218959
rect 48041 218931 48069 218959
rect 47979 218869 48007 218897
rect 48041 218869 48069 218897
rect 47979 218807 48007 218835
rect 48041 218807 48069 218835
rect 47979 218745 48007 218773
rect 48041 218745 48069 218773
rect 63339 218931 63367 218959
rect 63401 218931 63429 218959
rect 63339 218869 63367 218897
rect 63401 218869 63429 218897
rect 63339 218807 63367 218835
rect 63401 218807 63429 218835
rect 63339 218745 63367 218773
rect 63401 218745 63429 218773
rect 78699 218931 78727 218959
rect 78761 218931 78789 218959
rect 78699 218869 78727 218897
rect 78761 218869 78789 218897
rect 78699 218807 78727 218835
rect 78761 218807 78789 218835
rect 78699 218745 78727 218773
rect 78761 218745 78789 218773
rect 94059 218931 94087 218959
rect 94121 218931 94149 218959
rect 94059 218869 94087 218897
rect 94121 218869 94149 218897
rect 94059 218807 94087 218835
rect 94121 218807 94149 218835
rect 94059 218745 94087 218773
rect 94121 218745 94149 218773
rect 109419 218931 109447 218959
rect 109481 218931 109509 218959
rect 109419 218869 109447 218897
rect 109481 218869 109509 218897
rect 109419 218807 109447 218835
rect 109481 218807 109509 218835
rect 109419 218745 109447 218773
rect 109481 218745 109509 218773
rect 124779 218931 124807 218959
rect 124841 218931 124869 218959
rect 124779 218869 124807 218897
rect 124841 218869 124869 218897
rect 124779 218807 124807 218835
rect 124841 218807 124869 218835
rect 124779 218745 124807 218773
rect 124841 218745 124869 218773
rect 140139 218931 140167 218959
rect 140201 218931 140229 218959
rect 140139 218869 140167 218897
rect 140201 218869 140229 218897
rect 140139 218807 140167 218835
rect 140201 218807 140229 218835
rect 140139 218745 140167 218773
rect 140201 218745 140229 218773
rect 155499 218931 155527 218959
rect 155561 218931 155589 218959
rect 155499 218869 155527 218897
rect 155561 218869 155589 218897
rect 155499 218807 155527 218835
rect 155561 218807 155589 218835
rect 155499 218745 155527 218773
rect 155561 218745 155589 218773
rect 170859 218931 170887 218959
rect 170921 218931 170949 218959
rect 170859 218869 170887 218897
rect 170921 218869 170949 218897
rect 170859 218807 170887 218835
rect 170921 218807 170949 218835
rect 170859 218745 170887 218773
rect 170921 218745 170949 218773
rect 186219 218931 186247 218959
rect 186281 218931 186309 218959
rect 186219 218869 186247 218897
rect 186281 218869 186309 218897
rect 186219 218807 186247 218835
rect 186281 218807 186309 218835
rect 186219 218745 186247 218773
rect 186281 218745 186309 218773
rect 201579 218931 201607 218959
rect 201641 218931 201669 218959
rect 201579 218869 201607 218897
rect 201641 218869 201669 218897
rect 201579 218807 201607 218835
rect 201641 218807 201669 218835
rect 201579 218745 201607 218773
rect 201641 218745 201669 218773
rect 216939 218931 216967 218959
rect 217001 218931 217029 218959
rect 216939 218869 216967 218897
rect 217001 218869 217029 218897
rect 216939 218807 216967 218835
rect 217001 218807 217029 218835
rect 216939 218745 216967 218773
rect 217001 218745 217029 218773
rect 232299 218931 232327 218959
rect 232361 218931 232389 218959
rect 232299 218869 232327 218897
rect 232361 218869 232389 218897
rect 232299 218807 232327 218835
rect 232361 218807 232389 218835
rect 232299 218745 232327 218773
rect 232361 218745 232389 218773
rect 247659 218931 247687 218959
rect 247721 218931 247749 218959
rect 247659 218869 247687 218897
rect 247721 218869 247749 218897
rect 247659 218807 247687 218835
rect 247721 218807 247749 218835
rect 247659 218745 247687 218773
rect 247721 218745 247749 218773
rect 254577 218931 254605 218959
rect 254639 218931 254667 218959
rect 254701 218931 254729 218959
rect 254763 218931 254791 218959
rect 254577 218869 254605 218897
rect 254639 218869 254667 218897
rect 254701 218869 254729 218897
rect 254763 218869 254791 218897
rect 254577 218807 254605 218835
rect 254639 218807 254667 218835
rect 254701 218807 254729 218835
rect 254763 218807 254791 218835
rect 254577 218745 254605 218773
rect 254639 218745 254667 218773
rect 254701 218745 254729 218773
rect 254763 218745 254791 218773
rect 31437 212931 31465 212959
rect 31499 212931 31527 212959
rect 31561 212931 31589 212959
rect 31623 212931 31651 212959
rect 31437 212869 31465 212897
rect 31499 212869 31527 212897
rect 31561 212869 31589 212897
rect 31623 212869 31651 212897
rect 31437 212807 31465 212835
rect 31499 212807 31527 212835
rect 31561 212807 31589 212835
rect 31623 212807 31651 212835
rect 31437 212745 31465 212773
rect 31499 212745 31527 212773
rect 31561 212745 31589 212773
rect 31623 212745 31651 212773
rect 40299 212931 40327 212959
rect 40361 212931 40389 212959
rect 40299 212869 40327 212897
rect 40361 212869 40389 212897
rect 40299 212807 40327 212835
rect 40361 212807 40389 212835
rect 40299 212745 40327 212773
rect 40361 212745 40389 212773
rect 55659 212931 55687 212959
rect 55721 212931 55749 212959
rect 55659 212869 55687 212897
rect 55721 212869 55749 212897
rect 55659 212807 55687 212835
rect 55721 212807 55749 212835
rect 55659 212745 55687 212773
rect 55721 212745 55749 212773
rect 71019 212931 71047 212959
rect 71081 212931 71109 212959
rect 71019 212869 71047 212897
rect 71081 212869 71109 212897
rect 71019 212807 71047 212835
rect 71081 212807 71109 212835
rect 71019 212745 71047 212773
rect 71081 212745 71109 212773
rect 86379 212931 86407 212959
rect 86441 212931 86469 212959
rect 86379 212869 86407 212897
rect 86441 212869 86469 212897
rect 86379 212807 86407 212835
rect 86441 212807 86469 212835
rect 86379 212745 86407 212773
rect 86441 212745 86469 212773
rect 101739 212931 101767 212959
rect 101801 212931 101829 212959
rect 101739 212869 101767 212897
rect 101801 212869 101829 212897
rect 101739 212807 101767 212835
rect 101801 212807 101829 212835
rect 101739 212745 101767 212773
rect 101801 212745 101829 212773
rect 117099 212931 117127 212959
rect 117161 212931 117189 212959
rect 117099 212869 117127 212897
rect 117161 212869 117189 212897
rect 117099 212807 117127 212835
rect 117161 212807 117189 212835
rect 117099 212745 117127 212773
rect 117161 212745 117189 212773
rect 132459 212931 132487 212959
rect 132521 212931 132549 212959
rect 132459 212869 132487 212897
rect 132521 212869 132549 212897
rect 132459 212807 132487 212835
rect 132521 212807 132549 212835
rect 132459 212745 132487 212773
rect 132521 212745 132549 212773
rect 147819 212931 147847 212959
rect 147881 212931 147909 212959
rect 147819 212869 147847 212897
rect 147881 212869 147909 212897
rect 147819 212807 147847 212835
rect 147881 212807 147909 212835
rect 147819 212745 147847 212773
rect 147881 212745 147909 212773
rect 163179 212931 163207 212959
rect 163241 212931 163269 212959
rect 163179 212869 163207 212897
rect 163241 212869 163269 212897
rect 163179 212807 163207 212835
rect 163241 212807 163269 212835
rect 163179 212745 163207 212773
rect 163241 212745 163269 212773
rect 178539 212931 178567 212959
rect 178601 212931 178629 212959
rect 178539 212869 178567 212897
rect 178601 212869 178629 212897
rect 178539 212807 178567 212835
rect 178601 212807 178629 212835
rect 178539 212745 178567 212773
rect 178601 212745 178629 212773
rect 193899 212931 193927 212959
rect 193961 212931 193989 212959
rect 193899 212869 193927 212897
rect 193961 212869 193989 212897
rect 193899 212807 193927 212835
rect 193961 212807 193989 212835
rect 193899 212745 193927 212773
rect 193961 212745 193989 212773
rect 209259 212931 209287 212959
rect 209321 212931 209349 212959
rect 209259 212869 209287 212897
rect 209321 212869 209349 212897
rect 209259 212807 209287 212835
rect 209321 212807 209349 212835
rect 209259 212745 209287 212773
rect 209321 212745 209349 212773
rect 224619 212931 224647 212959
rect 224681 212931 224709 212959
rect 224619 212869 224647 212897
rect 224681 212869 224709 212897
rect 224619 212807 224647 212835
rect 224681 212807 224709 212835
rect 224619 212745 224647 212773
rect 224681 212745 224709 212773
rect 239979 212931 240007 212959
rect 240041 212931 240069 212959
rect 239979 212869 240007 212897
rect 240041 212869 240069 212897
rect 239979 212807 240007 212835
rect 240041 212807 240069 212835
rect 239979 212745 240007 212773
rect 240041 212745 240069 212773
rect 32619 209931 32647 209959
rect 32681 209931 32709 209959
rect 32619 209869 32647 209897
rect 32681 209869 32709 209897
rect 32619 209807 32647 209835
rect 32681 209807 32709 209835
rect 32619 209745 32647 209773
rect 32681 209745 32709 209773
rect 47979 209931 48007 209959
rect 48041 209931 48069 209959
rect 47979 209869 48007 209897
rect 48041 209869 48069 209897
rect 47979 209807 48007 209835
rect 48041 209807 48069 209835
rect 47979 209745 48007 209773
rect 48041 209745 48069 209773
rect 63339 209931 63367 209959
rect 63401 209931 63429 209959
rect 63339 209869 63367 209897
rect 63401 209869 63429 209897
rect 63339 209807 63367 209835
rect 63401 209807 63429 209835
rect 63339 209745 63367 209773
rect 63401 209745 63429 209773
rect 78699 209931 78727 209959
rect 78761 209931 78789 209959
rect 78699 209869 78727 209897
rect 78761 209869 78789 209897
rect 78699 209807 78727 209835
rect 78761 209807 78789 209835
rect 78699 209745 78727 209773
rect 78761 209745 78789 209773
rect 94059 209931 94087 209959
rect 94121 209931 94149 209959
rect 94059 209869 94087 209897
rect 94121 209869 94149 209897
rect 94059 209807 94087 209835
rect 94121 209807 94149 209835
rect 94059 209745 94087 209773
rect 94121 209745 94149 209773
rect 109419 209931 109447 209959
rect 109481 209931 109509 209959
rect 109419 209869 109447 209897
rect 109481 209869 109509 209897
rect 109419 209807 109447 209835
rect 109481 209807 109509 209835
rect 109419 209745 109447 209773
rect 109481 209745 109509 209773
rect 124779 209931 124807 209959
rect 124841 209931 124869 209959
rect 124779 209869 124807 209897
rect 124841 209869 124869 209897
rect 124779 209807 124807 209835
rect 124841 209807 124869 209835
rect 124779 209745 124807 209773
rect 124841 209745 124869 209773
rect 140139 209931 140167 209959
rect 140201 209931 140229 209959
rect 140139 209869 140167 209897
rect 140201 209869 140229 209897
rect 140139 209807 140167 209835
rect 140201 209807 140229 209835
rect 140139 209745 140167 209773
rect 140201 209745 140229 209773
rect 155499 209931 155527 209959
rect 155561 209931 155589 209959
rect 155499 209869 155527 209897
rect 155561 209869 155589 209897
rect 155499 209807 155527 209835
rect 155561 209807 155589 209835
rect 155499 209745 155527 209773
rect 155561 209745 155589 209773
rect 170859 209931 170887 209959
rect 170921 209931 170949 209959
rect 170859 209869 170887 209897
rect 170921 209869 170949 209897
rect 170859 209807 170887 209835
rect 170921 209807 170949 209835
rect 170859 209745 170887 209773
rect 170921 209745 170949 209773
rect 186219 209931 186247 209959
rect 186281 209931 186309 209959
rect 186219 209869 186247 209897
rect 186281 209869 186309 209897
rect 186219 209807 186247 209835
rect 186281 209807 186309 209835
rect 186219 209745 186247 209773
rect 186281 209745 186309 209773
rect 201579 209931 201607 209959
rect 201641 209931 201669 209959
rect 201579 209869 201607 209897
rect 201641 209869 201669 209897
rect 201579 209807 201607 209835
rect 201641 209807 201669 209835
rect 201579 209745 201607 209773
rect 201641 209745 201669 209773
rect 216939 209931 216967 209959
rect 217001 209931 217029 209959
rect 216939 209869 216967 209897
rect 217001 209869 217029 209897
rect 216939 209807 216967 209835
rect 217001 209807 217029 209835
rect 216939 209745 216967 209773
rect 217001 209745 217029 209773
rect 232299 209931 232327 209959
rect 232361 209931 232389 209959
rect 232299 209869 232327 209897
rect 232361 209869 232389 209897
rect 232299 209807 232327 209835
rect 232361 209807 232389 209835
rect 232299 209745 232327 209773
rect 232361 209745 232389 209773
rect 247659 209931 247687 209959
rect 247721 209931 247749 209959
rect 247659 209869 247687 209897
rect 247721 209869 247749 209897
rect 247659 209807 247687 209835
rect 247721 209807 247749 209835
rect 247659 209745 247687 209773
rect 247721 209745 247749 209773
rect 254577 209931 254605 209959
rect 254639 209931 254667 209959
rect 254701 209931 254729 209959
rect 254763 209931 254791 209959
rect 254577 209869 254605 209897
rect 254639 209869 254667 209897
rect 254701 209869 254729 209897
rect 254763 209869 254791 209897
rect 254577 209807 254605 209835
rect 254639 209807 254667 209835
rect 254701 209807 254729 209835
rect 254763 209807 254791 209835
rect 254577 209745 254605 209773
rect 254639 209745 254667 209773
rect 254701 209745 254729 209773
rect 254763 209745 254791 209773
rect 31437 203931 31465 203959
rect 31499 203931 31527 203959
rect 31561 203931 31589 203959
rect 31623 203931 31651 203959
rect 31437 203869 31465 203897
rect 31499 203869 31527 203897
rect 31561 203869 31589 203897
rect 31623 203869 31651 203897
rect 31437 203807 31465 203835
rect 31499 203807 31527 203835
rect 31561 203807 31589 203835
rect 31623 203807 31651 203835
rect 31437 203745 31465 203773
rect 31499 203745 31527 203773
rect 31561 203745 31589 203773
rect 31623 203745 31651 203773
rect 40299 203931 40327 203959
rect 40361 203931 40389 203959
rect 40299 203869 40327 203897
rect 40361 203869 40389 203897
rect 40299 203807 40327 203835
rect 40361 203807 40389 203835
rect 40299 203745 40327 203773
rect 40361 203745 40389 203773
rect 55659 203931 55687 203959
rect 55721 203931 55749 203959
rect 55659 203869 55687 203897
rect 55721 203869 55749 203897
rect 55659 203807 55687 203835
rect 55721 203807 55749 203835
rect 55659 203745 55687 203773
rect 55721 203745 55749 203773
rect 71019 203931 71047 203959
rect 71081 203931 71109 203959
rect 71019 203869 71047 203897
rect 71081 203869 71109 203897
rect 71019 203807 71047 203835
rect 71081 203807 71109 203835
rect 71019 203745 71047 203773
rect 71081 203745 71109 203773
rect 86379 203931 86407 203959
rect 86441 203931 86469 203959
rect 86379 203869 86407 203897
rect 86441 203869 86469 203897
rect 86379 203807 86407 203835
rect 86441 203807 86469 203835
rect 86379 203745 86407 203773
rect 86441 203745 86469 203773
rect 101739 203931 101767 203959
rect 101801 203931 101829 203959
rect 101739 203869 101767 203897
rect 101801 203869 101829 203897
rect 101739 203807 101767 203835
rect 101801 203807 101829 203835
rect 101739 203745 101767 203773
rect 101801 203745 101829 203773
rect 117099 203931 117127 203959
rect 117161 203931 117189 203959
rect 117099 203869 117127 203897
rect 117161 203869 117189 203897
rect 117099 203807 117127 203835
rect 117161 203807 117189 203835
rect 117099 203745 117127 203773
rect 117161 203745 117189 203773
rect 132459 203931 132487 203959
rect 132521 203931 132549 203959
rect 132459 203869 132487 203897
rect 132521 203869 132549 203897
rect 132459 203807 132487 203835
rect 132521 203807 132549 203835
rect 132459 203745 132487 203773
rect 132521 203745 132549 203773
rect 147819 203931 147847 203959
rect 147881 203931 147909 203959
rect 147819 203869 147847 203897
rect 147881 203869 147909 203897
rect 147819 203807 147847 203835
rect 147881 203807 147909 203835
rect 147819 203745 147847 203773
rect 147881 203745 147909 203773
rect 163179 203931 163207 203959
rect 163241 203931 163269 203959
rect 163179 203869 163207 203897
rect 163241 203869 163269 203897
rect 163179 203807 163207 203835
rect 163241 203807 163269 203835
rect 163179 203745 163207 203773
rect 163241 203745 163269 203773
rect 178539 203931 178567 203959
rect 178601 203931 178629 203959
rect 178539 203869 178567 203897
rect 178601 203869 178629 203897
rect 178539 203807 178567 203835
rect 178601 203807 178629 203835
rect 178539 203745 178567 203773
rect 178601 203745 178629 203773
rect 193899 203931 193927 203959
rect 193961 203931 193989 203959
rect 193899 203869 193927 203897
rect 193961 203869 193989 203897
rect 193899 203807 193927 203835
rect 193961 203807 193989 203835
rect 193899 203745 193927 203773
rect 193961 203745 193989 203773
rect 209259 203931 209287 203959
rect 209321 203931 209349 203959
rect 209259 203869 209287 203897
rect 209321 203869 209349 203897
rect 209259 203807 209287 203835
rect 209321 203807 209349 203835
rect 209259 203745 209287 203773
rect 209321 203745 209349 203773
rect 224619 203931 224647 203959
rect 224681 203931 224709 203959
rect 224619 203869 224647 203897
rect 224681 203869 224709 203897
rect 224619 203807 224647 203835
rect 224681 203807 224709 203835
rect 224619 203745 224647 203773
rect 224681 203745 224709 203773
rect 239979 203931 240007 203959
rect 240041 203931 240069 203959
rect 239979 203869 240007 203897
rect 240041 203869 240069 203897
rect 239979 203807 240007 203835
rect 240041 203807 240069 203835
rect 239979 203745 240007 203773
rect 240041 203745 240069 203773
rect 32619 200931 32647 200959
rect 32681 200931 32709 200959
rect 32619 200869 32647 200897
rect 32681 200869 32709 200897
rect 32619 200807 32647 200835
rect 32681 200807 32709 200835
rect 32619 200745 32647 200773
rect 32681 200745 32709 200773
rect 47979 200931 48007 200959
rect 48041 200931 48069 200959
rect 47979 200869 48007 200897
rect 48041 200869 48069 200897
rect 47979 200807 48007 200835
rect 48041 200807 48069 200835
rect 47979 200745 48007 200773
rect 48041 200745 48069 200773
rect 63339 200931 63367 200959
rect 63401 200931 63429 200959
rect 63339 200869 63367 200897
rect 63401 200869 63429 200897
rect 63339 200807 63367 200835
rect 63401 200807 63429 200835
rect 63339 200745 63367 200773
rect 63401 200745 63429 200773
rect 78699 200931 78727 200959
rect 78761 200931 78789 200959
rect 78699 200869 78727 200897
rect 78761 200869 78789 200897
rect 78699 200807 78727 200835
rect 78761 200807 78789 200835
rect 78699 200745 78727 200773
rect 78761 200745 78789 200773
rect 94059 200931 94087 200959
rect 94121 200931 94149 200959
rect 94059 200869 94087 200897
rect 94121 200869 94149 200897
rect 94059 200807 94087 200835
rect 94121 200807 94149 200835
rect 94059 200745 94087 200773
rect 94121 200745 94149 200773
rect 109419 200931 109447 200959
rect 109481 200931 109509 200959
rect 109419 200869 109447 200897
rect 109481 200869 109509 200897
rect 109419 200807 109447 200835
rect 109481 200807 109509 200835
rect 109419 200745 109447 200773
rect 109481 200745 109509 200773
rect 124779 200931 124807 200959
rect 124841 200931 124869 200959
rect 124779 200869 124807 200897
rect 124841 200869 124869 200897
rect 124779 200807 124807 200835
rect 124841 200807 124869 200835
rect 124779 200745 124807 200773
rect 124841 200745 124869 200773
rect 140139 200931 140167 200959
rect 140201 200931 140229 200959
rect 140139 200869 140167 200897
rect 140201 200869 140229 200897
rect 140139 200807 140167 200835
rect 140201 200807 140229 200835
rect 140139 200745 140167 200773
rect 140201 200745 140229 200773
rect 155499 200931 155527 200959
rect 155561 200931 155589 200959
rect 155499 200869 155527 200897
rect 155561 200869 155589 200897
rect 155499 200807 155527 200835
rect 155561 200807 155589 200835
rect 155499 200745 155527 200773
rect 155561 200745 155589 200773
rect 170859 200931 170887 200959
rect 170921 200931 170949 200959
rect 170859 200869 170887 200897
rect 170921 200869 170949 200897
rect 170859 200807 170887 200835
rect 170921 200807 170949 200835
rect 170859 200745 170887 200773
rect 170921 200745 170949 200773
rect 186219 200931 186247 200959
rect 186281 200931 186309 200959
rect 186219 200869 186247 200897
rect 186281 200869 186309 200897
rect 186219 200807 186247 200835
rect 186281 200807 186309 200835
rect 186219 200745 186247 200773
rect 186281 200745 186309 200773
rect 201579 200931 201607 200959
rect 201641 200931 201669 200959
rect 201579 200869 201607 200897
rect 201641 200869 201669 200897
rect 201579 200807 201607 200835
rect 201641 200807 201669 200835
rect 201579 200745 201607 200773
rect 201641 200745 201669 200773
rect 216939 200931 216967 200959
rect 217001 200931 217029 200959
rect 216939 200869 216967 200897
rect 217001 200869 217029 200897
rect 216939 200807 216967 200835
rect 217001 200807 217029 200835
rect 216939 200745 216967 200773
rect 217001 200745 217029 200773
rect 232299 200931 232327 200959
rect 232361 200931 232389 200959
rect 232299 200869 232327 200897
rect 232361 200869 232389 200897
rect 232299 200807 232327 200835
rect 232361 200807 232389 200835
rect 232299 200745 232327 200773
rect 232361 200745 232389 200773
rect 247659 200931 247687 200959
rect 247721 200931 247749 200959
rect 247659 200869 247687 200897
rect 247721 200869 247749 200897
rect 247659 200807 247687 200835
rect 247721 200807 247749 200835
rect 247659 200745 247687 200773
rect 247721 200745 247749 200773
rect 254577 200931 254605 200959
rect 254639 200931 254667 200959
rect 254701 200931 254729 200959
rect 254763 200931 254791 200959
rect 254577 200869 254605 200897
rect 254639 200869 254667 200897
rect 254701 200869 254729 200897
rect 254763 200869 254791 200897
rect 254577 200807 254605 200835
rect 254639 200807 254667 200835
rect 254701 200807 254729 200835
rect 254763 200807 254791 200835
rect 254577 200745 254605 200773
rect 254639 200745 254667 200773
rect 254701 200745 254729 200773
rect 254763 200745 254791 200773
rect 31437 194931 31465 194959
rect 31499 194931 31527 194959
rect 31561 194931 31589 194959
rect 31623 194931 31651 194959
rect 31437 194869 31465 194897
rect 31499 194869 31527 194897
rect 31561 194869 31589 194897
rect 31623 194869 31651 194897
rect 31437 194807 31465 194835
rect 31499 194807 31527 194835
rect 31561 194807 31589 194835
rect 31623 194807 31651 194835
rect 31437 194745 31465 194773
rect 31499 194745 31527 194773
rect 31561 194745 31589 194773
rect 31623 194745 31651 194773
rect 40299 194931 40327 194959
rect 40361 194931 40389 194959
rect 40299 194869 40327 194897
rect 40361 194869 40389 194897
rect 40299 194807 40327 194835
rect 40361 194807 40389 194835
rect 40299 194745 40327 194773
rect 40361 194745 40389 194773
rect 55659 194931 55687 194959
rect 55721 194931 55749 194959
rect 55659 194869 55687 194897
rect 55721 194869 55749 194897
rect 55659 194807 55687 194835
rect 55721 194807 55749 194835
rect 55659 194745 55687 194773
rect 55721 194745 55749 194773
rect 71019 194931 71047 194959
rect 71081 194931 71109 194959
rect 71019 194869 71047 194897
rect 71081 194869 71109 194897
rect 71019 194807 71047 194835
rect 71081 194807 71109 194835
rect 71019 194745 71047 194773
rect 71081 194745 71109 194773
rect 86379 194931 86407 194959
rect 86441 194931 86469 194959
rect 86379 194869 86407 194897
rect 86441 194869 86469 194897
rect 86379 194807 86407 194835
rect 86441 194807 86469 194835
rect 86379 194745 86407 194773
rect 86441 194745 86469 194773
rect 101739 194931 101767 194959
rect 101801 194931 101829 194959
rect 101739 194869 101767 194897
rect 101801 194869 101829 194897
rect 101739 194807 101767 194835
rect 101801 194807 101829 194835
rect 101739 194745 101767 194773
rect 101801 194745 101829 194773
rect 117099 194931 117127 194959
rect 117161 194931 117189 194959
rect 117099 194869 117127 194897
rect 117161 194869 117189 194897
rect 117099 194807 117127 194835
rect 117161 194807 117189 194835
rect 117099 194745 117127 194773
rect 117161 194745 117189 194773
rect 132459 194931 132487 194959
rect 132521 194931 132549 194959
rect 132459 194869 132487 194897
rect 132521 194869 132549 194897
rect 132459 194807 132487 194835
rect 132521 194807 132549 194835
rect 132459 194745 132487 194773
rect 132521 194745 132549 194773
rect 147819 194931 147847 194959
rect 147881 194931 147909 194959
rect 147819 194869 147847 194897
rect 147881 194869 147909 194897
rect 147819 194807 147847 194835
rect 147881 194807 147909 194835
rect 147819 194745 147847 194773
rect 147881 194745 147909 194773
rect 163179 194931 163207 194959
rect 163241 194931 163269 194959
rect 163179 194869 163207 194897
rect 163241 194869 163269 194897
rect 163179 194807 163207 194835
rect 163241 194807 163269 194835
rect 163179 194745 163207 194773
rect 163241 194745 163269 194773
rect 178539 194931 178567 194959
rect 178601 194931 178629 194959
rect 178539 194869 178567 194897
rect 178601 194869 178629 194897
rect 178539 194807 178567 194835
rect 178601 194807 178629 194835
rect 178539 194745 178567 194773
rect 178601 194745 178629 194773
rect 193899 194931 193927 194959
rect 193961 194931 193989 194959
rect 193899 194869 193927 194897
rect 193961 194869 193989 194897
rect 193899 194807 193927 194835
rect 193961 194807 193989 194835
rect 193899 194745 193927 194773
rect 193961 194745 193989 194773
rect 209259 194931 209287 194959
rect 209321 194931 209349 194959
rect 209259 194869 209287 194897
rect 209321 194869 209349 194897
rect 209259 194807 209287 194835
rect 209321 194807 209349 194835
rect 209259 194745 209287 194773
rect 209321 194745 209349 194773
rect 224619 194931 224647 194959
rect 224681 194931 224709 194959
rect 224619 194869 224647 194897
rect 224681 194869 224709 194897
rect 224619 194807 224647 194835
rect 224681 194807 224709 194835
rect 224619 194745 224647 194773
rect 224681 194745 224709 194773
rect 239979 194931 240007 194959
rect 240041 194931 240069 194959
rect 239979 194869 240007 194897
rect 240041 194869 240069 194897
rect 239979 194807 240007 194835
rect 240041 194807 240069 194835
rect 239979 194745 240007 194773
rect 240041 194745 240069 194773
rect 32619 191931 32647 191959
rect 32681 191931 32709 191959
rect 32619 191869 32647 191897
rect 32681 191869 32709 191897
rect 32619 191807 32647 191835
rect 32681 191807 32709 191835
rect 32619 191745 32647 191773
rect 32681 191745 32709 191773
rect 47979 191931 48007 191959
rect 48041 191931 48069 191959
rect 47979 191869 48007 191897
rect 48041 191869 48069 191897
rect 47979 191807 48007 191835
rect 48041 191807 48069 191835
rect 47979 191745 48007 191773
rect 48041 191745 48069 191773
rect 63339 191931 63367 191959
rect 63401 191931 63429 191959
rect 63339 191869 63367 191897
rect 63401 191869 63429 191897
rect 63339 191807 63367 191835
rect 63401 191807 63429 191835
rect 63339 191745 63367 191773
rect 63401 191745 63429 191773
rect 78699 191931 78727 191959
rect 78761 191931 78789 191959
rect 78699 191869 78727 191897
rect 78761 191869 78789 191897
rect 78699 191807 78727 191835
rect 78761 191807 78789 191835
rect 78699 191745 78727 191773
rect 78761 191745 78789 191773
rect 94059 191931 94087 191959
rect 94121 191931 94149 191959
rect 94059 191869 94087 191897
rect 94121 191869 94149 191897
rect 94059 191807 94087 191835
rect 94121 191807 94149 191835
rect 94059 191745 94087 191773
rect 94121 191745 94149 191773
rect 109419 191931 109447 191959
rect 109481 191931 109509 191959
rect 109419 191869 109447 191897
rect 109481 191869 109509 191897
rect 109419 191807 109447 191835
rect 109481 191807 109509 191835
rect 109419 191745 109447 191773
rect 109481 191745 109509 191773
rect 124779 191931 124807 191959
rect 124841 191931 124869 191959
rect 124779 191869 124807 191897
rect 124841 191869 124869 191897
rect 124779 191807 124807 191835
rect 124841 191807 124869 191835
rect 124779 191745 124807 191773
rect 124841 191745 124869 191773
rect 140139 191931 140167 191959
rect 140201 191931 140229 191959
rect 140139 191869 140167 191897
rect 140201 191869 140229 191897
rect 140139 191807 140167 191835
rect 140201 191807 140229 191835
rect 140139 191745 140167 191773
rect 140201 191745 140229 191773
rect 155499 191931 155527 191959
rect 155561 191931 155589 191959
rect 155499 191869 155527 191897
rect 155561 191869 155589 191897
rect 155499 191807 155527 191835
rect 155561 191807 155589 191835
rect 155499 191745 155527 191773
rect 155561 191745 155589 191773
rect 170859 191931 170887 191959
rect 170921 191931 170949 191959
rect 170859 191869 170887 191897
rect 170921 191869 170949 191897
rect 170859 191807 170887 191835
rect 170921 191807 170949 191835
rect 170859 191745 170887 191773
rect 170921 191745 170949 191773
rect 186219 191931 186247 191959
rect 186281 191931 186309 191959
rect 186219 191869 186247 191897
rect 186281 191869 186309 191897
rect 186219 191807 186247 191835
rect 186281 191807 186309 191835
rect 186219 191745 186247 191773
rect 186281 191745 186309 191773
rect 201579 191931 201607 191959
rect 201641 191931 201669 191959
rect 201579 191869 201607 191897
rect 201641 191869 201669 191897
rect 201579 191807 201607 191835
rect 201641 191807 201669 191835
rect 201579 191745 201607 191773
rect 201641 191745 201669 191773
rect 216939 191931 216967 191959
rect 217001 191931 217029 191959
rect 216939 191869 216967 191897
rect 217001 191869 217029 191897
rect 216939 191807 216967 191835
rect 217001 191807 217029 191835
rect 216939 191745 216967 191773
rect 217001 191745 217029 191773
rect 232299 191931 232327 191959
rect 232361 191931 232389 191959
rect 232299 191869 232327 191897
rect 232361 191869 232389 191897
rect 232299 191807 232327 191835
rect 232361 191807 232389 191835
rect 232299 191745 232327 191773
rect 232361 191745 232389 191773
rect 247659 191931 247687 191959
rect 247721 191931 247749 191959
rect 247659 191869 247687 191897
rect 247721 191869 247749 191897
rect 247659 191807 247687 191835
rect 247721 191807 247749 191835
rect 247659 191745 247687 191773
rect 247721 191745 247749 191773
rect 254577 191931 254605 191959
rect 254639 191931 254667 191959
rect 254701 191931 254729 191959
rect 254763 191931 254791 191959
rect 254577 191869 254605 191897
rect 254639 191869 254667 191897
rect 254701 191869 254729 191897
rect 254763 191869 254791 191897
rect 254577 191807 254605 191835
rect 254639 191807 254667 191835
rect 254701 191807 254729 191835
rect 254763 191807 254791 191835
rect 254577 191745 254605 191773
rect 254639 191745 254667 191773
rect 254701 191745 254729 191773
rect 254763 191745 254791 191773
rect 31437 185931 31465 185959
rect 31499 185931 31527 185959
rect 31561 185931 31589 185959
rect 31623 185931 31651 185959
rect 31437 185869 31465 185897
rect 31499 185869 31527 185897
rect 31561 185869 31589 185897
rect 31623 185869 31651 185897
rect 31437 185807 31465 185835
rect 31499 185807 31527 185835
rect 31561 185807 31589 185835
rect 31623 185807 31651 185835
rect 31437 185745 31465 185773
rect 31499 185745 31527 185773
rect 31561 185745 31589 185773
rect 31623 185745 31651 185773
rect 40299 185931 40327 185959
rect 40361 185931 40389 185959
rect 40299 185869 40327 185897
rect 40361 185869 40389 185897
rect 40299 185807 40327 185835
rect 40361 185807 40389 185835
rect 40299 185745 40327 185773
rect 40361 185745 40389 185773
rect 55659 185931 55687 185959
rect 55721 185931 55749 185959
rect 55659 185869 55687 185897
rect 55721 185869 55749 185897
rect 55659 185807 55687 185835
rect 55721 185807 55749 185835
rect 55659 185745 55687 185773
rect 55721 185745 55749 185773
rect 71019 185931 71047 185959
rect 71081 185931 71109 185959
rect 71019 185869 71047 185897
rect 71081 185869 71109 185897
rect 71019 185807 71047 185835
rect 71081 185807 71109 185835
rect 71019 185745 71047 185773
rect 71081 185745 71109 185773
rect 86379 185931 86407 185959
rect 86441 185931 86469 185959
rect 86379 185869 86407 185897
rect 86441 185869 86469 185897
rect 86379 185807 86407 185835
rect 86441 185807 86469 185835
rect 86379 185745 86407 185773
rect 86441 185745 86469 185773
rect 101739 185931 101767 185959
rect 101801 185931 101829 185959
rect 101739 185869 101767 185897
rect 101801 185869 101829 185897
rect 101739 185807 101767 185835
rect 101801 185807 101829 185835
rect 101739 185745 101767 185773
rect 101801 185745 101829 185773
rect 117099 185931 117127 185959
rect 117161 185931 117189 185959
rect 117099 185869 117127 185897
rect 117161 185869 117189 185897
rect 117099 185807 117127 185835
rect 117161 185807 117189 185835
rect 117099 185745 117127 185773
rect 117161 185745 117189 185773
rect 132459 185931 132487 185959
rect 132521 185931 132549 185959
rect 132459 185869 132487 185897
rect 132521 185869 132549 185897
rect 132459 185807 132487 185835
rect 132521 185807 132549 185835
rect 132459 185745 132487 185773
rect 132521 185745 132549 185773
rect 147819 185931 147847 185959
rect 147881 185931 147909 185959
rect 147819 185869 147847 185897
rect 147881 185869 147909 185897
rect 147819 185807 147847 185835
rect 147881 185807 147909 185835
rect 147819 185745 147847 185773
rect 147881 185745 147909 185773
rect 163179 185931 163207 185959
rect 163241 185931 163269 185959
rect 163179 185869 163207 185897
rect 163241 185869 163269 185897
rect 163179 185807 163207 185835
rect 163241 185807 163269 185835
rect 163179 185745 163207 185773
rect 163241 185745 163269 185773
rect 178539 185931 178567 185959
rect 178601 185931 178629 185959
rect 178539 185869 178567 185897
rect 178601 185869 178629 185897
rect 178539 185807 178567 185835
rect 178601 185807 178629 185835
rect 178539 185745 178567 185773
rect 178601 185745 178629 185773
rect 193899 185931 193927 185959
rect 193961 185931 193989 185959
rect 193899 185869 193927 185897
rect 193961 185869 193989 185897
rect 193899 185807 193927 185835
rect 193961 185807 193989 185835
rect 193899 185745 193927 185773
rect 193961 185745 193989 185773
rect 209259 185931 209287 185959
rect 209321 185931 209349 185959
rect 209259 185869 209287 185897
rect 209321 185869 209349 185897
rect 209259 185807 209287 185835
rect 209321 185807 209349 185835
rect 209259 185745 209287 185773
rect 209321 185745 209349 185773
rect 224619 185931 224647 185959
rect 224681 185931 224709 185959
rect 224619 185869 224647 185897
rect 224681 185869 224709 185897
rect 224619 185807 224647 185835
rect 224681 185807 224709 185835
rect 224619 185745 224647 185773
rect 224681 185745 224709 185773
rect 239979 185931 240007 185959
rect 240041 185931 240069 185959
rect 239979 185869 240007 185897
rect 240041 185869 240069 185897
rect 239979 185807 240007 185835
rect 240041 185807 240069 185835
rect 239979 185745 240007 185773
rect 240041 185745 240069 185773
rect 32619 182931 32647 182959
rect 32681 182931 32709 182959
rect 32619 182869 32647 182897
rect 32681 182869 32709 182897
rect 32619 182807 32647 182835
rect 32681 182807 32709 182835
rect 32619 182745 32647 182773
rect 32681 182745 32709 182773
rect 47979 182931 48007 182959
rect 48041 182931 48069 182959
rect 47979 182869 48007 182897
rect 48041 182869 48069 182897
rect 47979 182807 48007 182835
rect 48041 182807 48069 182835
rect 47979 182745 48007 182773
rect 48041 182745 48069 182773
rect 63339 182931 63367 182959
rect 63401 182931 63429 182959
rect 63339 182869 63367 182897
rect 63401 182869 63429 182897
rect 63339 182807 63367 182835
rect 63401 182807 63429 182835
rect 63339 182745 63367 182773
rect 63401 182745 63429 182773
rect 78699 182931 78727 182959
rect 78761 182931 78789 182959
rect 78699 182869 78727 182897
rect 78761 182869 78789 182897
rect 78699 182807 78727 182835
rect 78761 182807 78789 182835
rect 78699 182745 78727 182773
rect 78761 182745 78789 182773
rect 94059 182931 94087 182959
rect 94121 182931 94149 182959
rect 94059 182869 94087 182897
rect 94121 182869 94149 182897
rect 94059 182807 94087 182835
rect 94121 182807 94149 182835
rect 94059 182745 94087 182773
rect 94121 182745 94149 182773
rect 109419 182931 109447 182959
rect 109481 182931 109509 182959
rect 109419 182869 109447 182897
rect 109481 182869 109509 182897
rect 109419 182807 109447 182835
rect 109481 182807 109509 182835
rect 109419 182745 109447 182773
rect 109481 182745 109509 182773
rect 124779 182931 124807 182959
rect 124841 182931 124869 182959
rect 124779 182869 124807 182897
rect 124841 182869 124869 182897
rect 124779 182807 124807 182835
rect 124841 182807 124869 182835
rect 124779 182745 124807 182773
rect 124841 182745 124869 182773
rect 140139 182931 140167 182959
rect 140201 182931 140229 182959
rect 140139 182869 140167 182897
rect 140201 182869 140229 182897
rect 140139 182807 140167 182835
rect 140201 182807 140229 182835
rect 140139 182745 140167 182773
rect 140201 182745 140229 182773
rect 155499 182931 155527 182959
rect 155561 182931 155589 182959
rect 155499 182869 155527 182897
rect 155561 182869 155589 182897
rect 155499 182807 155527 182835
rect 155561 182807 155589 182835
rect 155499 182745 155527 182773
rect 155561 182745 155589 182773
rect 170859 182931 170887 182959
rect 170921 182931 170949 182959
rect 170859 182869 170887 182897
rect 170921 182869 170949 182897
rect 170859 182807 170887 182835
rect 170921 182807 170949 182835
rect 170859 182745 170887 182773
rect 170921 182745 170949 182773
rect 186219 182931 186247 182959
rect 186281 182931 186309 182959
rect 186219 182869 186247 182897
rect 186281 182869 186309 182897
rect 186219 182807 186247 182835
rect 186281 182807 186309 182835
rect 186219 182745 186247 182773
rect 186281 182745 186309 182773
rect 201579 182931 201607 182959
rect 201641 182931 201669 182959
rect 201579 182869 201607 182897
rect 201641 182869 201669 182897
rect 201579 182807 201607 182835
rect 201641 182807 201669 182835
rect 201579 182745 201607 182773
rect 201641 182745 201669 182773
rect 216939 182931 216967 182959
rect 217001 182931 217029 182959
rect 216939 182869 216967 182897
rect 217001 182869 217029 182897
rect 216939 182807 216967 182835
rect 217001 182807 217029 182835
rect 216939 182745 216967 182773
rect 217001 182745 217029 182773
rect 232299 182931 232327 182959
rect 232361 182931 232389 182959
rect 232299 182869 232327 182897
rect 232361 182869 232389 182897
rect 232299 182807 232327 182835
rect 232361 182807 232389 182835
rect 232299 182745 232327 182773
rect 232361 182745 232389 182773
rect 247659 182931 247687 182959
rect 247721 182931 247749 182959
rect 247659 182869 247687 182897
rect 247721 182869 247749 182897
rect 247659 182807 247687 182835
rect 247721 182807 247749 182835
rect 247659 182745 247687 182773
rect 247721 182745 247749 182773
rect 254577 182931 254605 182959
rect 254639 182931 254667 182959
rect 254701 182931 254729 182959
rect 254763 182931 254791 182959
rect 254577 182869 254605 182897
rect 254639 182869 254667 182897
rect 254701 182869 254729 182897
rect 254763 182869 254791 182897
rect 254577 182807 254605 182835
rect 254639 182807 254667 182835
rect 254701 182807 254729 182835
rect 254763 182807 254791 182835
rect 254577 182745 254605 182773
rect 254639 182745 254667 182773
rect 254701 182745 254729 182773
rect 254763 182745 254791 182773
rect 31437 176931 31465 176959
rect 31499 176931 31527 176959
rect 31561 176931 31589 176959
rect 31623 176931 31651 176959
rect 31437 176869 31465 176897
rect 31499 176869 31527 176897
rect 31561 176869 31589 176897
rect 31623 176869 31651 176897
rect 31437 176807 31465 176835
rect 31499 176807 31527 176835
rect 31561 176807 31589 176835
rect 31623 176807 31651 176835
rect 31437 176745 31465 176773
rect 31499 176745 31527 176773
rect 31561 176745 31589 176773
rect 31623 176745 31651 176773
rect 40299 176931 40327 176959
rect 40361 176931 40389 176959
rect 40299 176869 40327 176897
rect 40361 176869 40389 176897
rect 40299 176807 40327 176835
rect 40361 176807 40389 176835
rect 40299 176745 40327 176773
rect 40361 176745 40389 176773
rect 55659 176931 55687 176959
rect 55721 176931 55749 176959
rect 55659 176869 55687 176897
rect 55721 176869 55749 176897
rect 55659 176807 55687 176835
rect 55721 176807 55749 176835
rect 55659 176745 55687 176773
rect 55721 176745 55749 176773
rect 71019 176931 71047 176959
rect 71081 176931 71109 176959
rect 71019 176869 71047 176897
rect 71081 176869 71109 176897
rect 71019 176807 71047 176835
rect 71081 176807 71109 176835
rect 71019 176745 71047 176773
rect 71081 176745 71109 176773
rect 86379 176931 86407 176959
rect 86441 176931 86469 176959
rect 86379 176869 86407 176897
rect 86441 176869 86469 176897
rect 86379 176807 86407 176835
rect 86441 176807 86469 176835
rect 86379 176745 86407 176773
rect 86441 176745 86469 176773
rect 101739 176931 101767 176959
rect 101801 176931 101829 176959
rect 101739 176869 101767 176897
rect 101801 176869 101829 176897
rect 101739 176807 101767 176835
rect 101801 176807 101829 176835
rect 101739 176745 101767 176773
rect 101801 176745 101829 176773
rect 117099 176931 117127 176959
rect 117161 176931 117189 176959
rect 117099 176869 117127 176897
rect 117161 176869 117189 176897
rect 117099 176807 117127 176835
rect 117161 176807 117189 176835
rect 117099 176745 117127 176773
rect 117161 176745 117189 176773
rect 132459 176931 132487 176959
rect 132521 176931 132549 176959
rect 132459 176869 132487 176897
rect 132521 176869 132549 176897
rect 132459 176807 132487 176835
rect 132521 176807 132549 176835
rect 132459 176745 132487 176773
rect 132521 176745 132549 176773
rect 147819 176931 147847 176959
rect 147881 176931 147909 176959
rect 147819 176869 147847 176897
rect 147881 176869 147909 176897
rect 147819 176807 147847 176835
rect 147881 176807 147909 176835
rect 147819 176745 147847 176773
rect 147881 176745 147909 176773
rect 163179 176931 163207 176959
rect 163241 176931 163269 176959
rect 163179 176869 163207 176897
rect 163241 176869 163269 176897
rect 163179 176807 163207 176835
rect 163241 176807 163269 176835
rect 163179 176745 163207 176773
rect 163241 176745 163269 176773
rect 178539 176931 178567 176959
rect 178601 176931 178629 176959
rect 178539 176869 178567 176897
rect 178601 176869 178629 176897
rect 178539 176807 178567 176835
rect 178601 176807 178629 176835
rect 178539 176745 178567 176773
rect 178601 176745 178629 176773
rect 193899 176931 193927 176959
rect 193961 176931 193989 176959
rect 193899 176869 193927 176897
rect 193961 176869 193989 176897
rect 193899 176807 193927 176835
rect 193961 176807 193989 176835
rect 193899 176745 193927 176773
rect 193961 176745 193989 176773
rect 209259 176931 209287 176959
rect 209321 176931 209349 176959
rect 209259 176869 209287 176897
rect 209321 176869 209349 176897
rect 209259 176807 209287 176835
rect 209321 176807 209349 176835
rect 209259 176745 209287 176773
rect 209321 176745 209349 176773
rect 224619 176931 224647 176959
rect 224681 176931 224709 176959
rect 224619 176869 224647 176897
rect 224681 176869 224709 176897
rect 224619 176807 224647 176835
rect 224681 176807 224709 176835
rect 224619 176745 224647 176773
rect 224681 176745 224709 176773
rect 239979 176931 240007 176959
rect 240041 176931 240069 176959
rect 239979 176869 240007 176897
rect 240041 176869 240069 176897
rect 239979 176807 240007 176835
rect 240041 176807 240069 176835
rect 239979 176745 240007 176773
rect 240041 176745 240069 176773
rect 32619 173931 32647 173959
rect 32681 173931 32709 173959
rect 32619 173869 32647 173897
rect 32681 173869 32709 173897
rect 32619 173807 32647 173835
rect 32681 173807 32709 173835
rect 32619 173745 32647 173773
rect 32681 173745 32709 173773
rect 47979 173931 48007 173959
rect 48041 173931 48069 173959
rect 47979 173869 48007 173897
rect 48041 173869 48069 173897
rect 47979 173807 48007 173835
rect 48041 173807 48069 173835
rect 47979 173745 48007 173773
rect 48041 173745 48069 173773
rect 63339 173931 63367 173959
rect 63401 173931 63429 173959
rect 63339 173869 63367 173897
rect 63401 173869 63429 173897
rect 63339 173807 63367 173835
rect 63401 173807 63429 173835
rect 63339 173745 63367 173773
rect 63401 173745 63429 173773
rect 78699 173931 78727 173959
rect 78761 173931 78789 173959
rect 78699 173869 78727 173897
rect 78761 173869 78789 173897
rect 78699 173807 78727 173835
rect 78761 173807 78789 173835
rect 78699 173745 78727 173773
rect 78761 173745 78789 173773
rect 94059 173931 94087 173959
rect 94121 173931 94149 173959
rect 94059 173869 94087 173897
rect 94121 173869 94149 173897
rect 94059 173807 94087 173835
rect 94121 173807 94149 173835
rect 94059 173745 94087 173773
rect 94121 173745 94149 173773
rect 109419 173931 109447 173959
rect 109481 173931 109509 173959
rect 109419 173869 109447 173897
rect 109481 173869 109509 173897
rect 109419 173807 109447 173835
rect 109481 173807 109509 173835
rect 109419 173745 109447 173773
rect 109481 173745 109509 173773
rect 124779 173931 124807 173959
rect 124841 173931 124869 173959
rect 124779 173869 124807 173897
rect 124841 173869 124869 173897
rect 124779 173807 124807 173835
rect 124841 173807 124869 173835
rect 124779 173745 124807 173773
rect 124841 173745 124869 173773
rect 140139 173931 140167 173959
rect 140201 173931 140229 173959
rect 140139 173869 140167 173897
rect 140201 173869 140229 173897
rect 140139 173807 140167 173835
rect 140201 173807 140229 173835
rect 140139 173745 140167 173773
rect 140201 173745 140229 173773
rect 155499 173931 155527 173959
rect 155561 173931 155589 173959
rect 155499 173869 155527 173897
rect 155561 173869 155589 173897
rect 155499 173807 155527 173835
rect 155561 173807 155589 173835
rect 155499 173745 155527 173773
rect 155561 173745 155589 173773
rect 170859 173931 170887 173959
rect 170921 173931 170949 173959
rect 170859 173869 170887 173897
rect 170921 173869 170949 173897
rect 170859 173807 170887 173835
rect 170921 173807 170949 173835
rect 170859 173745 170887 173773
rect 170921 173745 170949 173773
rect 186219 173931 186247 173959
rect 186281 173931 186309 173959
rect 186219 173869 186247 173897
rect 186281 173869 186309 173897
rect 186219 173807 186247 173835
rect 186281 173807 186309 173835
rect 186219 173745 186247 173773
rect 186281 173745 186309 173773
rect 201579 173931 201607 173959
rect 201641 173931 201669 173959
rect 201579 173869 201607 173897
rect 201641 173869 201669 173897
rect 201579 173807 201607 173835
rect 201641 173807 201669 173835
rect 201579 173745 201607 173773
rect 201641 173745 201669 173773
rect 216939 173931 216967 173959
rect 217001 173931 217029 173959
rect 216939 173869 216967 173897
rect 217001 173869 217029 173897
rect 216939 173807 216967 173835
rect 217001 173807 217029 173835
rect 216939 173745 216967 173773
rect 217001 173745 217029 173773
rect 232299 173931 232327 173959
rect 232361 173931 232389 173959
rect 232299 173869 232327 173897
rect 232361 173869 232389 173897
rect 232299 173807 232327 173835
rect 232361 173807 232389 173835
rect 232299 173745 232327 173773
rect 232361 173745 232389 173773
rect 247659 173931 247687 173959
rect 247721 173931 247749 173959
rect 247659 173869 247687 173897
rect 247721 173869 247749 173897
rect 247659 173807 247687 173835
rect 247721 173807 247749 173835
rect 247659 173745 247687 173773
rect 247721 173745 247749 173773
rect 254577 173931 254605 173959
rect 254639 173931 254667 173959
rect 254701 173931 254729 173959
rect 254763 173931 254791 173959
rect 254577 173869 254605 173897
rect 254639 173869 254667 173897
rect 254701 173869 254729 173897
rect 254763 173869 254791 173897
rect 254577 173807 254605 173835
rect 254639 173807 254667 173835
rect 254701 173807 254729 173835
rect 254763 173807 254791 173835
rect 254577 173745 254605 173773
rect 254639 173745 254667 173773
rect 254701 173745 254729 173773
rect 254763 173745 254791 173773
rect 31437 167931 31465 167959
rect 31499 167931 31527 167959
rect 31561 167931 31589 167959
rect 31623 167931 31651 167959
rect 31437 167869 31465 167897
rect 31499 167869 31527 167897
rect 31561 167869 31589 167897
rect 31623 167869 31651 167897
rect 31437 167807 31465 167835
rect 31499 167807 31527 167835
rect 31561 167807 31589 167835
rect 31623 167807 31651 167835
rect 31437 167745 31465 167773
rect 31499 167745 31527 167773
rect 31561 167745 31589 167773
rect 31623 167745 31651 167773
rect 40299 167931 40327 167959
rect 40361 167931 40389 167959
rect 40299 167869 40327 167897
rect 40361 167869 40389 167897
rect 40299 167807 40327 167835
rect 40361 167807 40389 167835
rect 40299 167745 40327 167773
rect 40361 167745 40389 167773
rect 55659 167931 55687 167959
rect 55721 167931 55749 167959
rect 55659 167869 55687 167897
rect 55721 167869 55749 167897
rect 55659 167807 55687 167835
rect 55721 167807 55749 167835
rect 55659 167745 55687 167773
rect 55721 167745 55749 167773
rect 71019 167931 71047 167959
rect 71081 167931 71109 167959
rect 71019 167869 71047 167897
rect 71081 167869 71109 167897
rect 71019 167807 71047 167835
rect 71081 167807 71109 167835
rect 71019 167745 71047 167773
rect 71081 167745 71109 167773
rect 86379 167931 86407 167959
rect 86441 167931 86469 167959
rect 86379 167869 86407 167897
rect 86441 167869 86469 167897
rect 86379 167807 86407 167835
rect 86441 167807 86469 167835
rect 86379 167745 86407 167773
rect 86441 167745 86469 167773
rect 101739 167931 101767 167959
rect 101801 167931 101829 167959
rect 101739 167869 101767 167897
rect 101801 167869 101829 167897
rect 101739 167807 101767 167835
rect 101801 167807 101829 167835
rect 101739 167745 101767 167773
rect 101801 167745 101829 167773
rect 117099 167931 117127 167959
rect 117161 167931 117189 167959
rect 117099 167869 117127 167897
rect 117161 167869 117189 167897
rect 117099 167807 117127 167835
rect 117161 167807 117189 167835
rect 117099 167745 117127 167773
rect 117161 167745 117189 167773
rect 132459 167931 132487 167959
rect 132521 167931 132549 167959
rect 132459 167869 132487 167897
rect 132521 167869 132549 167897
rect 132459 167807 132487 167835
rect 132521 167807 132549 167835
rect 132459 167745 132487 167773
rect 132521 167745 132549 167773
rect 147819 167931 147847 167959
rect 147881 167931 147909 167959
rect 147819 167869 147847 167897
rect 147881 167869 147909 167897
rect 147819 167807 147847 167835
rect 147881 167807 147909 167835
rect 147819 167745 147847 167773
rect 147881 167745 147909 167773
rect 163179 167931 163207 167959
rect 163241 167931 163269 167959
rect 163179 167869 163207 167897
rect 163241 167869 163269 167897
rect 163179 167807 163207 167835
rect 163241 167807 163269 167835
rect 163179 167745 163207 167773
rect 163241 167745 163269 167773
rect 178539 167931 178567 167959
rect 178601 167931 178629 167959
rect 178539 167869 178567 167897
rect 178601 167869 178629 167897
rect 178539 167807 178567 167835
rect 178601 167807 178629 167835
rect 178539 167745 178567 167773
rect 178601 167745 178629 167773
rect 193899 167931 193927 167959
rect 193961 167931 193989 167959
rect 193899 167869 193927 167897
rect 193961 167869 193989 167897
rect 193899 167807 193927 167835
rect 193961 167807 193989 167835
rect 193899 167745 193927 167773
rect 193961 167745 193989 167773
rect 209259 167931 209287 167959
rect 209321 167931 209349 167959
rect 209259 167869 209287 167897
rect 209321 167869 209349 167897
rect 209259 167807 209287 167835
rect 209321 167807 209349 167835
rect 209259 167745 209287 167773
rect 209321 167745 209349 167773
rect 224619 167931 224647 167959
rect 224681 167931 224709 167959
rect 224619 167869 224647 167897
rect 224681 167869 224709 167897
rect 224619 167807 224647 167835
rect 224681 167807 224709 167835
rect 224619 167745 224647 167773
rect 224681 167745 224709 167773
rect 239979 167931 240007 167959
rect 240041 167931 240069 167959
rect 239979 167869 240007 167897
rect 240041 167869 240069 167897
rect 239979 167807 240007 167835
rect 240041 167807 240069 167835
rect 239979 167745 240007 167773
rect 240041 167745 240069 167773
rect 32619 164931 32647 164959
rect 32681 164931 32709 164959
rect 32619 164869 32647 164897
rect 32681 164869 32709 164897
rect 32619 164807 32647 164835
rect 32681 164807 32709 164835
rect 32619 164745 32647 164773
rect 32681 164745 32709 164773
rect 47979 164931 48007 164959
rect 48041 164931 48069 164959
rect 47979 164869 48007 164897
rect 48041 164869 48069 164897
rect 47979 164807 48007 164835
rect 48041 164807 48069 164835
rect 47979 164745 48007 164773
rect 48041 164745 48069 164773
rect 63339 164931 63367 164959
rect 63401 164931 63429 164959
rect 63339 164869 63367 164897
rect 63401 164869 63429 164897
rect 63339 164807 63367 164835
rect 63401 164807 63429 164835
rect 63339 164745 63367 164773
rect 63401 164745 63429 164773
rect 78699 164931 78727 164959
rect 78761 164931 78789 164959
rect 78699 164869 78727 164897
rect 78761 164869 78789 164897
rect 78699 164807 78727 164835
rect 78761 164807 78789 164835
rect 78699 164745 78727 164773
rect 78761 164745 78789 164773
rect 94059 164931 94087 164959
rect 94121 164931 94149 164959
rect 94059 164869 94087 164897
rect 94121 164869 94149 164897
rect 94059 164807 94087 164835
rect 94121 164807 94149 164835
rect 94059 164745 94087 164773
rect 94121 164745 94149 164773
rect 109419 164931 109447 164959
rect 109481 164931 109509 164959
rect 109419 164869 109447 164897
rect 109481 164869 109509 164897
rect 109419 164807 109447 164835
rect 109481 164807 109509 164835
rect 109419 164745 109447 164773
rect 109481 164745 109509 164773
rect 124779 164931 124807 164959
rect 124841 164931 124869 164959
rect 124779 164869 124807 164897
rect 124841 164869 124869 164897
rect 124779 164807 124807 164835
rect 124841 164807 124869 164835
rect 124779 164745 124807 164773
rect 124841 164745 124869 164773
rect 140139 164931 140167 164959
rect 140201 164931 140229 164959
rect 140139 164869 140167 164897
rect 140201 164869 140229 164897
rect 140139 164807 140167 164835
rect 140201 164807 140229 164835
rect 140139 164745 140167 164773
rect 140201 164745 140229 164773
rect 155499 164931 155527 164959
rect 155561 164931 155589 164959
rect 155499 164869 155527 164897
rect 155561 164869 155589 164897
rect 155499 164807 155527 164835
rect 155561 164807 155589 164835
rect 155499 164745 155527 164773
rect 155561 164745 155589 164773
rect 170859 164931 170887 164959
rect 170921 164931 170949 164959
rect 170859 164869 170887 164897
rect 170921 164869 170949 164897
rect 170859 164807 170887 164835
rect 170921 164807 170949 164835
rect 170859 164745 170887 164773
rect 170921 164745 170949 164773
rect 186219 164931 186247 164959
rect 186281 164931 186309 164959
rect 186219 164869 186247 164897
rect 186281 164869 186309 164897
rect 186219 164807 186247 164835
rect 186281 164807 186309 164835
rect 186219 164745 186247 164773
rect 186281 164745 186309 164773
rect 201579 164931 201607 164959
rect 201641 164931 201669 164959
rect 201579 164869 201607 164897
rect 201641 164869 201669 164897
rect 201579 164807 201607 164835
rect 201641 164807 201669 164835
rect 201579 164745 201607 164773
rect 201641 164745 201669 164773
rect 216939 164931 216967 164959
rect 217001 164931 217029 164959
rect 216939 164869 216967 164897
rect 217001 164869 217029 164897
rect 216939 164807 216967 164835
rect 217001 164807 217029 164835
rect 216939 164745 216967 164773
rect 217001 164745 217029 164773
rect 232299 164931 232327 164959
rect 232361 164931 232389 164959
rect 232299 164869 232327 164897
rect 232361 164869 232389 164897
rect 232299 164807 232327 164835
rect 232361 164807 232389 164835
rect 232299 164745 232327 164773
rect 232361 164745 232389 164773
rect 247659 164931 247687 164959
rect 247721 164931 247749 164959
rect 247659 164869 247687 164897
rect 247721 164869 247749 164897
rect 247659 164807 247687 164835
rect 247721 164807 247749 164835
rect 247659 164745 247687 164773
rect 247721 164745 247749 164773
rect 254577 164931 254605 164959
rect 254639 164931 254667 164959
rect 254701 164931 254729 164959
rect 254763 164931 254791 164959
rect 254577 164869 254605 164897
rect 254639 164869 254667 164897
rect 254701 164869 254729 164897
rect 254763 164869 254791 164897
rect 254577 164807 254605 164835
rect 254639 164807 254667 164835
rect 254701 164807 254729 164835
rect 254763 164807 254791 164835
rect 254577 164745 254605 164773
rect 254639 164745 254667 164773
rect 254701 164745 254729 164773
rect 254763 164745 254791 164773
rect 31437 158931 31465 158959
rect 31499 158931 31527 158959
rect 31561 158931 31589 158959
rect 31623 158931 31651 158959
rect 31437 158869 31465 158897
rect 31499 158869 31527 158897
rect 31561 158869 31589 158897
rect 31623 158869 31651 158897
rect 31437 158807 31465 158835
rect 31499 158807 31527 158835
rect 31561 158807 31589 158835
rect 31623 158807 31651 158835
rect 31437 158745 31465 158773
rect 31499 158745 31527 158773
rect 31561 158745 31589 158773
rect 31623 158745 31651 158773
rect 40299 158931 40327 158959
rect 40361 158931 40389 158959
rect 40299 158869 40327 158897
rect 40361 158869 40389 158897
rect 40299 158807 40327 158835
rect 40361 158807 40389 158835
rect 40299 158745 40327 158773
rect 40361 158745 40389 158773
rect 55659 158931 55687 158959
rect 55721 158931 55749 158959
rect 55659 158869 55687 158897
rect 55721 158869 55749 158897
rect 55659 158807 55687 158835
rect 55721 158807 55749 158835
rect 55659 158745 55687 158773
rect 55721 158745 55749 158773
rect 71019 158931 71047 158959
rect 71081 158931 71109 158959
rect 71019 158869 71047 158897
rect 71081 158869 71109 158897
rect 71019 158807 71047 158835
rect 71081 158807 71109 158835
rect 71019 158745 71047 158773
rect 71081 158745 71109 158773
rect 86379 158931 86407 158959
rect 86441 158931 86469 158959
rect 86379 158869 86407 158897
rect 86441 158869 86469 158897
rect 86379 158807 86407 158835
rect 86441 158807 86469 158835
rect 86379 158745 86407 158773
rect 86441 158745 86469 158773
rect 101739 158931 101767 158959
rect 101801 158931 101829 158959
rect 101739 158869 101767 158897
rect 101801 158869 101829 158897
rect 101739 158807 101767 158835
rect 101801 158807 101829 158835
rect 101739 158745 101767 158773
rect 101801 158745 101829 158773
rect 117099 158931 117127 158959
rect 117161 158931 117189 158959
rect 117099 158869 117127 158897
rect 117161 158869 117189 158897
rect 117099 158807 117127 158835
rect 117161 158807 117189 158835
rect 117099 158745 117127 158773
rect 117161 158745 117189 158773
rect 132459 158931 132487 158959
rect 132521 158931 132549 158959
rect 132459 158869 132487 158897
rect 132521 158869 132549 158897
rect 132459 158807 132487 158835
rect 132521 158807 132549 158835
rect 132459 158745 132487 158773
rect 132521 158745 132549 158773
rect 147819 158931 147847 158959
rect 147881 158931 147909 158959
rect 147819 158869 147847 158897
rect 147881 158869 147909 158897
rect 147819 158807 147847 158835
rect 147881 158807 147909 158835
rect 147819 158745 147847 158773
rect 147881 158745 147909 158773
rect 163179 158931 163207 158959
rect 163241 158931 163269 158959
rect 163179 158869 163207 158897
rect 163241 158869 163269 158897
rect 163179 158807 163207 158835
rect 163241 158807 163269 158835
rect 163179 158745 163207 158773
rect 163241 158745 163269 158773
rect 178539 158931 178567 158959
rect 178601 158931 178629 158959
rect 178539 158869 178567 158897
rect 178601 158869 178629 158897
rect 178539 158807 178567 158835
rect 178601 158807 178629 158835
rect 178539 158745 178567 158773
rect 178601 158745 178629 158773
rect 193899 158931 193927 158959
rect 193961 158931 193989 158959
rect 193899 158869 193927 158897
rect 193961 158869 193989 158897
rect 193899 158807 193927 158835
rect 193961 158807 193989 158835
rect 193899 158745 193927 158773
rect 193961 158745 193989 158773
rect 209259 158931 209287 158959
rect 209321 158931 209349 158959
rect 209259 158869 209287 158897
rect 209321 158869 209349 158897
rect 209259 158807 209287 158835
rect 209321 158807 209349 158835
rect 209259 158745 209287 158773
rect 209321 158745 209349 158773
rect 224619 158931 224647 158959
rect 224681 158931 224709 158959
rect 224619 158869 224647 158897
rect 224681 158869 224709 158897
rect 224619 158807 224647 158835
rect 224681 158807 224709 158835
rect 224619 158745 224647 158773
rect 224681 158745 224709 158773
rect 239979 158931 240007 158959
rect 240041 158931 240069 158959
rect 239979 158869 240007 158897
rect 240041 158869 240069 158897
rect 239979 158807 240007 158835
rect 240041 158807 240069 158835
rect 239979 158745 240007 158773
rect 240041 158745 240069 158773
rect 32619 155931 32647 155959
rect 32681 155931 32709 155959
rect 32619 155869 32647 155897
rect 32681 155869 32709 155897
rect 32619 155807 32647 155835
rect 32681 155807 32709 155835
rect 32619 155745 32647 155773
rect 32681 155745 32709 155773
rect 47979 155931 48007 155959
rect 48041 155931 48069 155959
rect 47979 155869 48007 155897
rect 48041 155869 48069 155897
rect 47979 155807 48007 155835
rect 48041 155807 48069 155835
rect 47979 155745 48007 155773
rect 48041 155745 48069 155773
rect 63339 155931 63367 155959
rect 63401 155931 63429 155959
rect 63339 155869 63367 155897
rect 63401 155869 63429 155897
rect 63339 155807 63367 155835
rect 63401 155807 63429 155835
rect 63339 155745 63367 155773
rect 63401 155745 63429 155773
rect 78699 155931 78727 155959
rect 78761 155931 78789 155959
rect 78699 155869 78727 155897
rect 78761 155869 78789 155897
rect 78699 155807 78727 155835
rect 78761 155807 78789 155835
rect 78699 155745 78727 155773
rect 78761 155745 78789 155773
rect 94059 155931 94087 155959
rect 94121 155931 94149 155959
rect 94059 155869 94087 155897
rect 94121 155869 94149 155897
rect 94059 155807 94087 155835
rect 94121 155807 94149 155835
rect 94059 155745 94087 155773
rect 94121 155745 94149 155773
rect 109419 155931 109447 155959
rect 109481 155931 109509 155959
rect 109419 155869 109447 155897
rect 109481 155869 109509 155897
rect 109419 155807 109447 155835
rect 109481 155807 109509 155835
rect 109419 155745 109447 155773
rect 109481 155745 109509 155773
rect 124779 155931 124807 155959
rect 124841 155931 124869 155959
rect 124779 155869 124807 155897
rect 124841 155869 124869 155897
rect 124779 155807 124807 155835
rect 124841 155807 124869 155835
rect 124779 155745 124807 155773
rect 124841 155745 124869 155773
rect 140139 155931 140167 155959
rect 140201 155931 140229 155959
rect 140139 155869 140167 155897
rect 140201 155869 140229 155897
rect 140139 155807 140167 155835
rect 140201 155807 140229 155835
rect 140139 155745 140167 155773
rect 140201 155745 140229 155773
rect 155499 155931 155527 155959
rect 155561 155931 155589 155959
rect 155499 155869 155527 155897
rect 155561 155869 155589 155897
rect 155499 155807 155527 155835
rect 155561 155807 155589 155835
rect 155499 155745 155527 155773
rect 155561 155745 155589 155773
rect 170859 155931 170887 155959
rect 170921 155931 170949 155959
rect 170859 155869 170887 155897
rect 170921 155869 170949 155897
rect 170859 155807 170887 155835
rect 170921 155807 170949 155835
rect 170859 155745 170887 155773
rect 170921 155745 170949 155773
rect 186219 155931 186247 155959
rect 186281 155931 186309 155959
rect 186219 155869 186247 155897
rect 186281 155869 186309 155897
rect 186219 155807 186247 155835
rect 186281 155807 186309 155835
rect 186219 155745 186247 155773
rect 186281 155745 186309 155773
rect 201579 155931 201607 155959
rect 201641 155931 201669 155959
rect 201579 155869 201607 155897
rect 201641 155869 201669 155897
rect 201579 155807 201607 155835
rect 201641 155807 201669 155835
rect 201579 155745 201607 155773
rect 201641 155745 201669 155773
rect 216939 155931 216967 155959
rect 217001 155931 217029 155959
rect 216939 155869 216967 155897
rect 217001 155869 217029 155897
rect 216939 155807 216967 155835
rect 217001 155807 217029 155835
rect 216939 155745 216967 155773
rect 217001 155745 217029 155773
rect 232299 155931 232327 155959
rect 232361 155931 232389 155959
rect 232299 155869 232327 155897
rect 232361 155869 232389 155897
rect 232299 155807 232327 155835
rect 232361 155807 232389 155835
rect 232299 155745 232327 155773
rect 232361 155745 232389 155773
rect 247659 155931 247687 155959
rect 247721 155931 247749 155959
rect 247659 155869 247687 155897
rect 247721 155869 247749 155897
rect 247659 155807 247687 155835
rect 247721 155807 247749 155835
rect 247659 155745 247687 155773
rect 247721 155745 247749 155773
rect 254577 155931 254605 155959
rect 254639 155931 254667 155959
rect 254701 155931 254729 155959
rect 254763 155931 254791 155959
rect 254577 155869 254605 155897
rect 254639 155869 254667 155897
rect 254701 155869 254729 155897
rect 254763 155869 254791 155897
rect 254577 155807 254605 155835
rect 254639 155807 254667 155835
rect 254701 155807 254729 155835
rect 254763 155807 254791 155835
rect 254577 155745 254605 155773
rect 254639 155745 254667 155773
rect 254701 155745 254729 155773
rect 254763 155745 254791 155773
rect 31437 149931 31465 149959
rect 31499 149931 31527 149959
rect 31561 149931 31589 149959
rect 31623 149931 31651 149959
rect 31437 149869 31465 149897
rect 31499 149869 31527 149897
rect 31561 149869 31589 149897
rect 31623 149869 31651 149897
rect 31437 149807 31465 149835
rect 31499 149807 31527 149835
rect 31561 149807 31589 149835
rect 31623 149807 31651 149835
rect 31437 149745 31465 149773
rect 31499 149745 31527 149773
rect 31561 149745 31589 149773
rect 31623 149745 31651 149773
rect 40299 149931 40327 149959
rect 40361 149931 40389 149959
rect 40299 149869 40327 149897
rect 40361 149869 40389 149897
rect 40299 149807 40327 149835
rect 40361 149807 40389 149835
rect 40299 149745 40327 149773
rect 40361 149745 40389 149773
rect 55659 149931 55687 149959
rect 55721 149931 55749 149959
rect 55659 149869 55687 149897
rect 55721 149869 55749 149897
rect 55659 149807 55687 149835
rect 55721 149807 55749 149835
rect 55659 149745 55687 149773
rect 55721 149745 55749 149773
rect 71019 149931 71047 149959
rect 71081 149931 71109 149959
rect 71019 149869 71047 149897
rect 71081 149869 71109 149897
rect 71019 149807 71047 149835
rect 71081 149807 71109 149835
rect 71019 149745 71047 149773
rect 71081 149745 71109 149773
rect 86379 149931 86407 149959
rect 86441 149931 86469 149959
rect 86379 149869 86407 149897
rect 86441 149869 86469 149897
rect 86379 149807 86407 149835
rect 86441 149807 86469 149835
rect 86379 149745 86407 149773
rect 86441 149745 86469 149773
rect 101739 149931 101767 149959
rect 101801 149931 101829 149959
rect 101739 149869 101767 149897
rect 101801 149869 101829 149897
rect 101739 149807 101767 149835
rect 101801 149807 101829 149835
rect 101739 149745 101767 149773
rect 101801 149745 101829 149773
rect 117099 149931 117127 149959
rect 117161 149931 117189 149959
rect 117099 149869 117127 149897
rect 117161 149869 117189 149897
rect 117099 149807 117127 149835
rect 117161 149807 117189 149835
rect 117099 149745 117127 149773
rect 117161 149745 117189 149773
rect 132459 149931 132487 149959
rect 132521 149931 132549 149959
rect 132459 149869 132487 149897
rect 132521 149869 132549 149897
rect 132459 149807 132487 149835
rect 132521 149807 132549 149835
rect 132459 149745 132487 149773
rect 132521 149745 132549 149773
rect 147819 149931 147847 149959
rect 147881 149931 147909 149959
rect 147819 149869 147847 149897
rect 147881 149869 147909 149897
rect 147819 149807 147847 149835
rect 147881 149807 147909 149835
rect 147819 149745 147847 149773
rect 147881 149745 147909 149773
rect 163179 149931 163207 149959
rect 163241 149931 163269 149959
rect 163179 149869 163207 149897
rect 163241 149869 163269 149897
rect 163179 149807 163207 149835
rect 163241 149807 163269 149835
rect 163179 149745 163207 149773
rect 163241 149745 163269 149773
rect 178539 149931 178567 149959
rect 178601 149931 178629 149959
rect 178539 149869 178567 149897
rect 178601 149869 178629 149897
rect 178539 149807 178567 149835
rect 178601 149807 178629 149835
rect 178539 149745 178567 149773
rect 178601 149745 178629 149773
rect 193899 149931 193927 149959
rect 193961 149931 193989 149959
rect 193899 149869 193927 149897
rect 193961 149869 193989 149897
rect 193899 149807 193927 149835
rect 193961 149807 193989 149835
rect 193899 149745 193927 149773
rect 193961 149745 193989 149773
rect 209259 149931 209287 149959
rect 209321 149931 209349 149959
rect 209259 149869 209287 149897
rect 209321 149869 209349 149897
rect 209259 149807 209287 149835
rect 209321 149807 209349 149835
rect 209259 149745 209287 149773
rect 209321 149745 209349 149773
rect 224619 149931 224647 149959
rect 224681 149931 224709 149959
rect 224619 149869 224647 149897
rect 224681 149869 224709 149897
rect 224619 149807 224647 149835
rect 224681 149807 224709 149835
rect 224619 149745 224647 149773
rect 224681 149745 224709 149773
rect 239979 149931 240007 149959
rect 240041 149931 240069 149959
rect 239979 149869 240007 149897
rect 240041 149869 240069 149897
rect 239979 149807 240007 149835
rect 240041 149807 240069 149835
rect 239979 149745 240007 149773
rect 240041 149745 240069 149773
rect 32619 146931 32647 146959
rect 32681 146931 32709 146959
rect 32619 146869 32647 146897
rect 32681 146869 32709 146897
rect 32619 146807 32647 146835
rect 32681 146807 32709 146835
rect 32619 146745 32647 146773
rect 32681 146745 32709 146773
rect 47979 146931 48007 146959
rect 48041 146931 48069 146959
rect 47979 146869 48007 146897
rect 48041 146869 48069 146897
rect 47979 146807 48007 146835
rect 48041 146807 48069 146835
rect 47979 146745 48007 146773
rect 48041 146745 48069 146773
rect 63339 146931 63367 146959
rect 63401 146931 63429 146959
rect 63339 146869 63367 146897
rect 63401 146869 63429 146897
rect 63339 146807 63367 146835
rect 63401 146807 63429 146835
rect 63339 146745 63367 146773
rect 63401 146745 63429 146773
rect 78699 146931 78727 146959
rect 78761 146931 78789 146959
rect 78699 146869 78727 146897
rect 78761 146869 78789 146897
rect 78699 146807 78727 146835
rect 78761 146807 78789 146835
rect 78699 146745 78727 146773
rect 78761 146745 78789 146773
rect 94059 146931 94087 146959
rect 94121 146931 94149 146959
rect 94059 146869 94087 146897
rect 94121 146869 94149 146897
rect 94059 146807 94087 146835
rect 94121 146807 94149 146835
rect 94059 146745 94087 146773
rect 94121 146745 94149 146773
rect 109419 146931 109447 146959
rect 109481 146931 109509 146959
rect 109419 146869 109447 146897
rect 109481 146869 109509 146897
rect 109419 146807 109447 146835
rect 109481 146807 109509 146835
rect 109419 146745 109447 146773
rect 109481 146745 109509 146773
rect 124779 146931 124807 146959
rect 124841 146931 124869 146959
rect 124779 146869 124807 146897
rect 124841 146869 124869 146897
rect 124779 146807 124807 146835
rect 124841 146807 124869 146835
rect 124779 146745 124807 146773
rect 124841 146745 124869 146773
rect 140139 146931 140167 146959
rect 140201 146931 140229 146959
rect 140139 146869 140167 146897
rect 140201 146869 140229 146897
rect 140139 146807 140167 146835
rect 140201 146807 140229 146835
rect 140139 146745 140167 146773
rect 140201 146745 140229 146773
rect 155499 146931 155527 146959
rect 155561 146931 155589 146959
rect 155499 146869 155527 146897
rect 155561 146869 155589 146897
rect 155499 146807 155527 146835
rect 155561 146807 155589 146835
rect 155499 146745 155527 146773
rect 155561 146745 155589 146773
rect 170859 146931 170887 146959
rect 170921 146931 170949 146959
rect 170859 146869 170887 146897
rect 170921 146869 170949 146897
rect 170859 146807 170887 146835
rect 170921 146807 170949 146835
rect 170859 146745 170887 146773
rect 170921 146745 170949 146773
rect 186219 146931 186247 146959
rect 186281 146931 186309 146959
rect 186219 146869 186247 146897
rect 186281 146869 186309 146897
rect 186219 146807 186247 146835
rect 186281 146807 186309 146835
rect 186219 146745 186247 146773
rect 186281 146745 186309 146773
rect 201579 146931 201607 146959
rect 201641 146931 201669 146959
rect 201579 146869 201607 146897
rect 201641 146869 201669 146897
rect 201579 146807 201607 146835
rect 201641 146807 201669 146835
rect 201579 146745 201607 146773
rect 201641 146745 201669 146773
rect 216939 146931 216967 146959
rect 217001 146931 217029 146959
rect 216939 146869 216967 146897
rect 217001 146869 217029 146897
rect 216939 146807 216967 146835
rect 217001 146807 217029 146835
rect 216939 146745 216967 146773
rect 217001 146745 217029 146773
rect 232299 146931 232327 146959
rect 232361 146931 232389 146959
rect 232299 146869 232327 146897
rect 232361 146869 232389 146897
rect 232299 146807 232327 146835
rect 232361 146807 232389 146835
rect 232299 146745 232327 146773
rect 232361 146745 232389 146773
rect 247659 146931 247687 146959
rect 247721 146931 247749 146959
rect 247659 146869 247687 146897
rect 247721 146869 247749 146897
rect 247659 146807 247687 146835
rect 247721 146807 247749 146835
rect 247659 146745 247687 146773
rect 247721 146745 247749 146773
rect 254577 146931 254605 146959
rect 254639 146931 254667 146959
rect 254701 146931 254729 146959
rect 254763 146931 254791 146959
rect 254577 146869 254605 146897
rect 254639 146869 254667 146897
rect 254701 146869 254729 146897
rect 254763 146869 254791 146897
rect 254577 146807 254605 146835
rect 254639 146807 254667 146835
rect 254701 146807 254729 146835
rect 254763 146807 254791 146835
rect 254577 146745 254605 146773
rect 254639 146745 254667 146773
rect 254701 146745 254729 146773
rect 254763 146745 254791 146773
rect 31437 140931 31465 140959
rect 31499 140931 31527 140959
rect 31561 140931 31589 140959
rect 31623 140931 31651 140959
rect 31437 140869 31465 140897
rect 31499 140869 31527 140897
rect 31561 140869 31589 140897
rect 31623 140869 31651 140897
rect 31437 140807 31465 140835
rect 31499 140807 31527 140835
rect 31561 140807 31589 140835
rect 31623 140807 31651 140835
rect 31437 140745 31465 140773
rect 31499 140745 31527 140773
rect 31561 140745 31589 140773
rect 31623 140745 31651 140773
rect 40299 140931 40327 140959
rect 40361 140931 40389 140959
rect 40299 140869 40327 140897
rect 40361 140869 40389 140897
rect 40299 140807 40327 140835
rect 40361 140807 40389 140835
rect 40299 140745 40327 140773
rect 40361 140745 40389 140773
rect 55659 140931 55687 140959
rect 55721 140931 55749 140959
rect 55659 140869 55687 140897
rect 55721 140869 55749 140897
rect 55659 140807 55687 140835
rect 55721 140807 55749 140835
rect 55659 140745 55687 140773
rect 55721 140745 55749 140773
rect 71019 140931 71047 140959
rect 71081 140931 71109 140959
rect 71019 140869 71047 140897
rect 71081 140869 71109 140897
rect 71019 140807 71047 140835
rect 71081 140807 71109 140835
rect 71019 140745 71047 140773
rect 71081 140745 71109 140773
rect 86379 140931 86407 140959
rect 86441 140931 86469 140959
rect 86379 140869 86407 140897
rect 86441 140869 86469 140897
rect 86379 140807 86407 140835
rect 86441 140807 86469 140835
rect 86379 140745 86407 140773
rect 86441 140745 86469 140773
rect 101739 140931 101767 140959
rect 101801 140931 101829 140959
rect 101739 140869 101767 140897
rect 101801 140869 101829 140897
rect 101739 140807 101767 140835
rect 101801 140807 101829 140835
rect 101739 140745 101767 140773
rect 101801 140745 101829 140773
rect 117099 140931 117127 140959
rect 117161 140931 117189 140959
rect 117099 140869 117127 140897
rect 117161 140869 117189 140897
rect 117099 140807 117127 140835
rect 117161 140807 117189 140835
rect 117099 140745 117127 140773
rect 117161 140745 117189 140773
rect 132459 140931 132487 140959
rect 132521 140931 132549 140959
rect 132459 140869 132487 140897
rect 132521 140869 132549 140897
rect 132459 140807 132487 140835
rect 132521 140807 132549 140835
rect 132459 140745 132487 140773
rect 132521 140745 132549 140773
rect 147819 140931 147847 140959
rect 147881 140931 147909 140959
rect 147819 140869 147847 140897
rect 147881 140869 147909 140897
rect 147819 140807 147847 140835
rect 147881 140807 147909 140835
rect 147819 140745 147847 140773
rect 147881 140745 147909 140773
rect 163179 140931 163207 140959
rect 163241 140931 163269 140959
rect 163179 140869 163207 140897
rect 163241 140869 163269 140897
rect 163179 140807 163207 140835
rect 163241 140807 163269 140835
rect 163179 140745 163207 140773
rect 163241 140745 163269 140773
rect 178539 140931 178567 140959
rect 178601 140931 178629 140959
rect 178539 140869 178567 140897
rect 178601 140869 178629 140897
rect 178539 140807 178567 140835
rect 178601 140807 178629 140835
rect 178539 140745 178567 140773
rect 178601 140745 178629 140773
rect 193899 140931 193927 140959
rect 193961 140931 193989 140959
rect 193899 140869 193927 140897
rect 193961 140869 193989 140897
rect 193899 140807 193927 140835
rect 193961 140807 193989 140835
rect 193899 140745 193927 140773
rect 193961 140745 193989 140773
rect 209259 140931 209287 140959
rect 209321 140931 209349 140959
rect 209259 140869 209287 140897
rect 209321 140869 209349 140897
rect 209259 140807 209287 140835
rect 209321 140807 209349 140835
rect 209259 140745 209287 140773
rect 209321 140745 209349 140773
rect 224619 140931 224647 140959
rect 224681 140931 224709 140959
rect 224619 140869 224647 140897
rect 224681 140869 224709 140897
rect 224619 140807 224647 140835
rect 224681 140807 224709 140835
rect 224619 140745 224647 140773
rect 224681 140745 224709 140773
rect 239979 140931 240007 140959
rect 240041 140931 240069 140959
rect 239979 140869 240007 140897
rect 240041 140869 240069 140897
rect 239979 140807 240007 140835
rect 240041 140807 240069 140835
rect 239979 140745 240007 140773
rect 240041 140745 240069 140773
rect 32619 137931 32647 137959
rect 32681 137931 32709 137959
rect 32619 137869 32647 137897
rect 32681 137869 32709 137897
rect 32619 137807 32647 137835
rect 32681 137807 32709 137835
rect 32619 137745 32647 137773
rect 32681 137745 32709 137773
rect 47979 137931 48007 137959
rect 48041 137931 48069 137959
rect 47979 137869 48007 137897
rect 48041 137869 48069 137897
rect 47979 137807 48007 137835
rect 48041 137807 48069 137835
rect 47979 137745 48007 137773
rect 48041 137745 48069 137773
rect 63339 137931 63367 137959
rect 63401 137931 63429 137959
rect 63339 137869 63367 137897
rect 63401 137869 63429 137897
rect 63339 137807 63367 137835
rect 63401 137807 63429 137835
rect 63339 137745 63367 137773
rect 63401 137745 63429 137773
rect 78699 137931 78727 137959
rect 78761 137931 78789 137959
rect 78699 137869 78727 137897
rect 78761 137869 78789 137897
rect 78699 137807 78727 137835
rect 78761 137807 78789 137835
rect 78699 137745 78727 137773
rect 78761 137745 78789 137773
rect 94059 137931 94087 137959
rect 94121 137931 94149 137959
rect 94059 137869 94087 137897
rect 94121 137869 94149 137897
rect 94059 137807 94087 137835
rect 94121 137807 94149 137835
rect 94059 137745 94087 137773
rect 94121 137745 94149 137773
rect 109419 137931 109447 137959
rect 109481 137931 109509 137959
rect 109419 137869 109447 137897
rect 109481 137869 109509 137897
rect 109419 137807 109447 137835
rect 109481 137807 109509 137835
rect 109419 137745 109447 137773
rect 109481 137745 109509 137773
rect 124779 137931 124807 137959
rect 124841 137931 124869 137959
rect 124779 137869 124807 137897
rect 124841 137869 124869 137897
rect 124779 137807 124807 137835
rect 124841 137807 124869 137835
rect 124779 137745 124807 137773
rect 124841 137745 124869 137773
rect 140139 137931 140167 137959
rect 140201 137931 140229 137959
rect 140139 137869 140167 137897
rect 140201 137869 140229 137897
rect 140139 137807 140167 137835
rect 140201 137807 140229 137835
rect 140139 137745 140167 137773
rect 140201 137745 140229 137773
rect 155499 137931 155527 137959
rect 155561 137931 155589 137959
rect 155499 137869 155527 137897
rect 155561 137869 155589 137897
rect 155499 137807 155527 137835
rect 155561 137807 155589 137835
rect 155499 137745 155527 137773
rect 155561 137745 155589 137773
rect 170859 137931 170887 137959
rect 170921 137931 170949 137959
rect 170859 137869 170887 137897
rect 170921 137869 170949 137897
rect 170859 137807 170887 137835
rect 170921 137807 170949 137835
rect 170859 137745 170887 137773
rect 170921 137745 170949 137773
rect 186219 137931 186247 137959
rect 186281 137931 186309 137959
rect 186219 137869 186247 137897
rect 186281 137869 186309 137897
rect 186219 137807 186247 137835
rect 186281 137807 186309 137835
rect 186219 137745 186247 137773
rect 186281 137745 186309 137773
rect 201579 137931 201607 137959
rect 201641 137931 201669 137959
rect 201579 137869 201607 137897
rect 201641 137869 201669 137897
rect 201579 137807 201607 137835
rect 201641 137807 201669 137835
rect 201579 137745 201607 137773
rect 201641 137745 201669 137773
rect 216939 137931 216967 137959
rect 217001 137931 217029 137959
rect 216939 137869 216967 137897
rect 217001 137869 217029 137897
rect 216939 137807 216967 137835
rect 217001 137807 217029 137835
rect 216939 137745 216967 137773
rect 217001 137745 217029 137773
rect 232299 137931 232327 137959
rect 232361 137931 232389 137959
rect 232299 137869 232327 137897
rect 232361 137869 232389 137897
rect 232299 137807 232327 137835
rect 232361 137807 232389 137835
rect 232299 137745 232327 137773
rect 232361 137745 232389 137773
rect 247659 137931 247687 137959
rect 247721 137931 247749 137959
rect 247659 137869 247687 137897
rect 247721 137869 247749 137897
rect 247659 137807 247687 137835
rect 247721 137807 247749 137835
rect 247659 137745 247687 137773
rect 247721 137745 247749 137773
rect 254577 137931 254605 137959
rect 254639 137931 254667 137959
rect 254701 137931 254729 137959
rect 254763 137931 254791 137959
rect 254577 137869 254605 137897
rect 254639 137869 254667 137897
rect 254701 137869 254729 137897
rect 254763 137869 254791 137897
rect 254577 137807 254605 137835
rect 254639 137807 254667 137835
rect 254701 137807 254729 137835
rect 254763 137807 254791 137835
rect 254577 137745 254605 137773
rect 254639 137745 254667 137773
rect 254701 137745 254729 137773
rect 254763 137745 254791 137773
rect 31437 131931 31465 131959
rect 31499 131931 31527 131959
rect 31561 131931 31589 131959
rect 31623 131931 31651 131959
rect 31437 131869 31465 131897
rect 31499 131869 31527 131897
rect 31561 131869 31589 131897
rect 31623 131869 31651 131897
rect 31437 131807 31465 131835
rect 31499 131807 31527 131835
rect 31561 131807 31589 131835
rect 31623 131807 31651 131835
rect 31437 131745 31465 131773
rect 31499 131745 31527 131773
rect 31561 131745 31589 131773
rect 31623 131745 31651 131773
rect 40299 131931 40327 131959
rect 40361 131931 40389 131959
rect 40299 131869 40327 131897
rect 40361 131869 40389 131897
rect 40299 131807 40327 131835
rect 40361 131807 40389 131835
rect 40299 131745 40327 131773
rect 40361 131745 40389 131773
rect 55659 131931 55687 131959
rect 55721 131931 55749 131959
rect 55659 131869 55687 131897
rect 55721 131869 55749 131897
rect 55659 131807 55687 131835
rect 55721 131807 55749 131835
rect 55659 131745 55687 131773
rect 55721 131745 55749 131773
rect 71019 131931 71047 131959
rect 71081 131931 71109 131959
rect 71019 131869 71047 131897
rect 71081 131869 71109 131897
rect 71019 131807 71047 131835
rect 71081 131807 71109 131835
rect 71019 131745 71047 131773
rect 71081 131745 71109 131773
rect 86379 131931 86407 131959
rect 86441 131931 86469 131959
rect 86379 131869 86407 131897
rect 86441 131869 86469 131897
rect 86379 131807 86407 131835
rect 86441 131807 86469 131835
rect 86379 131745 86407 131773
rect 86441 131745 86469 131773
rect 101739 131931 101767 131959
rect 101801 131931 101829 131959
rect 101739 131869 101767 131897
rect 101801 131869 101829 131897
rect 101739 131807 101767 131835
rect 101801 131807 101829 131835
rect 101739 131745 101767 131773
rect 101801 131745 101829 131773
rect 117099 131931 117127 131959
rect 117161 131931 117189 131959
rect 117099 131869 117127 131897
rect 117161 131869 117189 131897
rect 117099 131807 117127 131835
rect 117161 131807 117189 131835
rect 117099 131745 117127 131773
rect 117161 131745 117189 131773
rect 132459 131931 132487 131959
rect 132521 131931 132549 131959
rect 132459 131869 132487 131897
rect 132521 131869 132549 131897
rect 132459 131807 132487 131835
rect 132521 131807 132549 131835
rect 132459 131745 132487 131773
rect 132521 131745 132549 131773
rect 147819 131931 147847 131959
rect 147881 131931 147909 131959
rect 147819 131869 147847 131897
rect 147881 131869 147909 131897
rect 147819 131807 147847 131835
rect 147881 131807 147909 131835
rect 147819 131745 147847 131773
rect 147881 131745 147909 131773
rect 163179 131931 163207 131959
rect 163241 131931 163269 131959
rect 163179 131869 163207 131897
rect 163241 131869 163269 131897
rect 163179 131807 163207 131835
rect 163241 131807 163269 131835
rect 163179 131745 163207 131773
rect 163241 131745 163269 131773
rect 178539 131931 178567 131959
rect 178601 131931 178629 131959
rect 178539 131869 178567 131897
rect 178601 131869 178629 131897
rect 178539 131807 178567 131835
rect 178601 131807 178629 131835
rect 178539 131745 178567 131773
rect 178601 131745 178629 131773
rect 193899 131931 193927 131959
rect 193961 131931 193989 131959
rect 193899 131869 193927 131897
rect 193961 131869 193989 131897
rect 193899 131807 193927 131835
rect 193961 131807 193989 131835
rect 193899 131745 193927 131773
rect 193961 131745 193989 131773
rect 209259 131931 209287 131959
rect 209321 131931 209349 131959
rect 209259 131869 209287 131897
rect 209321 131869 209349 131897
rect 209259 131807 209287 131835
rect 209321 131807 209349 131835
rect 209259 131745 209287 131773
rect 209321 131745 209349 131773
rect 224619 131931 224647 131959
rect 224681 131931 224709 131959
rect 224619 131869 224647 131897
rect 224681 131869 224709 131897
rect 224619 131807 224647 131835
rect 224681 131807 224709 131835
rect 224619 131745 224647 131773
rect 224681 131745 224709 131773
rect 239979 131931 240007 131959
rect 240041 131931 240069 131959
rect 239979 131869 240007 131897
rect 240041 131869 240069 131897
rect 239979 131807 240007 131835
rect 240041 131807 240069 131835
rect 239979 131745 240007 131773
rect 240041 131745 240069 131773
rect 32619 128931 32647 128959
rect 32681 128931 32709 128959
rect 32619 128869 32647 128897
rect 32681 128869 32709 128897
rect 32619 128807 32647 128835
rect 32681 128807 32709 128835
rect 32619 128745 32647 128773
rect 32681 128745 32709 128773
rect 47979 128931 48007 128959
rect 48041 128931 48069 128959
rect 47979 128869 48007 128897
rect 48041 128869 48069 128897
rect 47979 128807 48007 128835
rect 48041 128807 48069 128835
rect 47979 128745 48007 128773
rect 48041 128745 48069 128773
rect 63339 128931 63367 128959
rect 63401 128931 63429 128959
rect 63339 128869 63367 128897
rect 63401 128869 63429 128897
rect 63339 128807 63367 128835
rect 63401 128807 63429 128835
rect 63339 128745 63367 128773
rect 63401 128745 63429 128773
rect 78699 128931 78727 128959
rect 78761 128931 78789 128959
rect 78699 128869 78727 128897
rect 78761 128869 78789 128897
rect 78699 128807 78727 128835
rect 78761 128807 78789 128835
rect 78699 128745 78727 128773
rect 78761 128745 78789 128773
rect 94059 128931 94087 128959
rect 94121 128931 94149 128959
rect 94059 128869 94087 128897
rect 94121 128869 94149 128897
rect 94059 128807 94087 128835
rect 94121 128807 94149 128835
rect 94059 128745 94087 128773
rect 94121 128745 94149 128773
rect 109419 128931 109447 128959
rect 109481 128931 109509 128959
rect 109419 128869 109447 128897
rect 109481 128869 109509 128897
rect 109419 128807 109447 128835
rect 109481 128807 109509 128835
rect 109419 128745 109447 128773
rect 109481 128745 109509 128773
rect 124779 128931 124807 128959
rect 124841 128931 124869 128959
rect 124779 128869 124807 128897
rect 124841 128869 124869 128897
rect 124779 128807 124807 128835
rect 124841 128807 124869 128835
rect 124779 128745 124807 128773
rect 124841 128745 124869 128773
rect 140139 128931 140167 128959
rect 140201 128931 140229 128959
rect 140139 128869 140167 128897
rect 140201 128869 140229 128897
rect 140139 128807 140167 128835
rect 140201 128807 140229 128835
rect 140139 128745 140167 128773
rect 140201 128745 140229 128773
rect 155499 128931 155527 128959
rect 155561 128931 155589 128959
rect 155499 128869 155527 128897
rect 155561 128869 155589 128897
rect 155499 128807 155527 128835
rect 155561 128807 155589 128835
rect 155499 128745 155527 128773
rect 155561 128745 155589 128773
rect 170859 128931 170887 128959
rect 170921 128931 170949 128959
rect 170859 128869 170887 128897
rect 170921 128869 170949 128897
rect 170859 128807 170887 128835
rect 170921 128807 170949 128835
rect 170859 128745 170887 128773
rect 170921 128745 170949 128773
rect 186219 128931 186247 128959
rect 186281 128931 186309 128959
rect 186219 128869 186247 128897
rect 186281 128869 186309 128897
rect 186219 128807 186247 128835
rect 186281 128807 186309 128835
rect 186219 128745 186247 128773
rect 186281 128745 186309 128773
rect 201579 128931 201607 128959
rect 201641 128931 201669 128959
rect 201579 128869 201607 128897
rect 201641 128869 201669 128897
rect 201579 128807 201607 128835
rect 201641 128807 201669 128835
rect 201579 128745 201607 128773
rect 201641 128745 201669 128773
rect 216939 128931 216967 128959
rect 217001 128931 217029 128959
rect 216939 128869 216967 128897
rect 217001 128869 217029 128897
rect 216939 128807 216967 128835
rect 217001 128807 217029 128835
rect 216939 128745 216967 128773
rect 217001 128745 217029 128773
rect 232299 128931 232327 128959
rect 232361 128931 232389 128959
rect 232299 128869 232327 128897
rect 232361 128869 232389 128897
rect 232299 128807 232327 128835
rect 232361 128807 232389 128835
rect 232299 128745 232327 128773
rect 232361 128745 232389 128773
rect 247659 128931 247687 128959
rect 247721 128931 247749 128959
rect 247659 128869 247687 128897
rect 247721 128869 247749 128897
rect 247659 128807 247687 128835
rect 247721 128807 247749 128835
rect 247659 128745 247687 128773
rect 247721 128745 247749 128773
rect 254577 128931 254605 128959
rect 254639 128931 254667 128959
rect 254701 128931 254729 128959
rect 254763 128931 254791 128959
rect 254577 128869 254605 128897
rect 254639 128869 254667 128897
rect 254701 128869 254729 128897
rect 254763 128869 254791 128897
rect 254577 128807 254605 128835
rect 254639 128807 254667 128835
rect 254701 128807 254729 128835
rect 254763 128807 254791 128835
rect 254577 128745 254605 128773
rect 254639 128745 254667 128773
rect 254701 128745 254729 128773
rect 254763 128745 254791 128773
rect 31437 122931 31465 122959
rect 31499 122931 31527 122959
rect 31561 122931 31589 122959
rect 31623 122931 31651 122959
rect 31437 122869 31465 122897
rect 31499 122869 31527 122897
rect 31561 122869 31589 122897
rect 31623 122869 31651 122897
rect 31437 122807 31465 122835
rect 31499 122807 31527 122835
rect 31561 122807 31589 122835
rect 31623 122807 31651 122835
rect 31437 122745 31465 122773
rect 31499 122745 31527 122773
rect 31561 122745 31589 122773
rect 31623 122745 31651 122773
rect 40299 122931 40327 122959
rect 40361 122931 40389 122959
rect 40299 122869 40327 122897
rect 40361 122869 40389 122897
rect 40299 122807 40327 122835
rect 40361 122807 40389 122835
rect 40299 122745 40327 122773
rect 40361 122745 40389 122773
rect 55659 122931 55687 122959
rect 55721 122931 55749 122959
rect 55659 122869 55687 122897
rect 55721 122869 55749 122897
rect 55659 122807 55687 122835
rect 55721 122807 55749 122835
rect 55659 122745 55687 122773
rect 55721 122745 55749 122773
rect 71019 122931 71047 122959
rect 71081 122931 71109 122959
rect 71019 122869 71047 122897
rect 71081 122869 71109 122897
rect 71019 122807 71047 122835
rect 71081 122807 71109 122835
rect 71019 122745 71047 122773
rect 71081 122745 71109 122773
rect 86379 122931 86407 122959
rect 86441 122931 86469 122959
rect 86379 122869 86407 122897
rect 86441 122869 86469 122897
rect 86379 122807 86407 122835
rect 86441 122807 86469 122835
rect 86379 122745 86407 122773
rect 86441 122745 86469 122773
rect 101739 122931 101767 122959
rect 101801 122931 101829 122959
rect 101739 122869 101767 122897
rect 101801 122869 101829 122897
rect 101739 122807 101767 122835
rect 101801 122807 101829 122835
rect 101739 122745 101767 122773
rect 101801 122745 101829 122773
rect 117099 122931 117127 122959
rect 117161 122931 117189 122959
rect 117099 122869 117127 122897
rect 117161 122869 117189 122897
rect 117099 122807 117127 122835
rect 117161 122807 117189 122835
rect 117099 122745 117127 122773
rect 117161 122745 117189 122773
rect 132459 122931 132487 122959
rect 132521 122931 132549 122959
rect 132459 122869 132487 122897
rect 132521 122869 132549 122897
rect 132459 122807 132487 122835
rect 132521 122807 132549 122835
rect 132459 122745 132487 122773
rect 132521 122745 132549 122773
rect 147819 122931 147847 122959
rect 147881 122931 147909 122959
rect 147819 122869 147847 122897
rect 147881 122869 147909 122897
rect 147819 122807 147847 122835
rect 147881 122807 147909 122835
rect 147819 122745 147847 122773
rect 147881 122745 147909 122773
rect 163179 122931 163207 122959
rect 163241 122931 163269 122959
rect 163179 122869 163207 122897
rect 163241 122869 163269 122897
rect 163179 122807 163207 122835
rect 163241 122807 163269 122835
rect 163179 122745 163207 122773
rect 163241 122745 163269 122773
rect 178539 122931 178567 122959
rect 178601 122931 178629 122959
rect 178539 122869 178567 122897
rect 178601 122869 178629 122897
rect 178539 122807 178567 122835
rect 178601 122807 178629 122835
rect 178539 122745 178567 122773
rect 178601 122745 178629 122773
rect 193899 122931 193927 122959
rect 193961 122931 193989 122959
rect 193899 122869 193927 122897
rect 193961 122869 193989 122897
rect 193899 122807 193927 122835
rect 193961 122807 193989 122835
rect 193899 122745 193927 122773
rect 193961 122745 193989 122773
rect 209259 122931 209287 122959
rect 209321 122931 209349 122959
rect 209259 122869 209287 122897
rect 209321 122869 209349 122897
rect 209259 122807 209287 122835
rect 209321 122807 209349 122835
rect 209259 122745 209287 122773
rect 209321 122745 209349 122773
rect 224619 122931 224647 122959
rect 224681 122931 224709 122959
rect 224619 122869 224647 122897
rect 224681 122869 224709 122897
rect 224619 122807 224647 122835
rect 224681 122807 224709 122835
rect 224619 122745 224647 122773
rect 224681 122745 224709 122773
rect 239979 122931 240007 122959
rect 240041 122931 240069 122959
rect 239979 122869 240007 122897
rect 240041 122869 240069 122897
rect 239979 122807 240007 122835
rect 240041 122807 240069 122835
rect 239979 122745 240007 122773
rect 240041 122745 240069 122773
rect 32619 119931 32647 119959
rect 32681 119931 32709 119959
rect 32619 119869 32647 119897
rect 32681 119869 32709 119897
rect 32619 119807 32647 119835
rect 32681 119807 32709 119835
rect 32619 119745 32647 119773
rect 32681 119745 32709 119773
rect 47979 119931 48007 119959
rect 48041 119931 48069 119959
rect 47979 119869 48007 119897
rect 48041 119869 48069 119897
rect 47979 119807 48007 119835
rect 48041 119807 48069 119835
rect 47979 119745 48007 119773
rect 48041 119745 48069 119773
rect 63339 119931 63367 119959
rect 63401 119931 63429 119959
rect 63339 119869 63367 119897
rect 63401 119869 63429 119897
rect 63339 119807 63367 119835
rect 63401 119807 63429 119835
rect 63339 119745 63367 119773
rect 63401 119745 63429 119773
rect 78699 119931 78727 119959
rect 78761 119931 78789 119959
rect 78699 119869 78727 119897
rect 78761 119869 78789 119897
rect 78699 119807 78727 119835
rect 78761 119807 78789 119835
rect 78699 119745 78727 119773
rect 78761 119745 78789 119773
rect 94059 119931 94087 119959
rect 94121 119931 94149 119959
rect 94059 119869 94087 119897
rect 94121 119869 94149 119897
rect 94059 119807 94087 119835
rect 94121 119807 94149 119835
rect 94059 119745 94087 119773
rect 94121 119745 94149 119773
rect 109419 119931 109447 119959
rect 109481 119931 109509 119959
rect 109419 119869 109447 119897
rect 109481 119869 109509 119897
rect 109419 119807 109447 119835
rect 109481 119807 109509 119835
rect 109419 119745 109447 119773
rect 109481 119745 109509 119773
rect 124779 119931 124807 119959
rect 124841 119931 124869 119959
rect 124779 119869 124807 119897
rect 124841 119869 124869 119897
rect 124779 119807 124807 119835
rect 124841 119807 124869 119835
rect 124779 119745 124807 119773
rect 124841 119745 124869 119773
rect 140139 119931 140167 119959
rect 140201 119931 140229 119959
rect 140139 119869 140167 119897
rect 140201 119869 140229 119897
rect 140139 119807 140167 119835
rect 140201 119807 140229 119835
rect 140139 119745 140167 119773
rect 140201 119745 140229 119773
rect 155499 119931 155527 119959
rect 155561 119931 155589 119959
rect 155499 119869 155527 119897
rect 155561 119869 155589 119897
rect 155499 119807 155527 119835
rect 155561 119807 155589 119835
rect 155499 119745 155527 119773
rect 155561 119745 155589 119773
rect 170859 119931 170887 119959
rect 170921 119931 170949 119959
rect 170859 119869 170887 119897
rect 170921 119869 170949 119897
rect 170859 119807 170887 119835
rect 170921 119807 170949 119835
rect 170859 119745 170887 119773
rect 170921 119745 170949 119773
rect 186219 119931 186247 119959
rect 186281 119931 186309 119959
rect 186219 119869 186247 119897
rect 186281 119869 186309 119897
rect 186219 119807 186247 119835
rect 186281 119807 186309 119835
rect 186219 119745 186247 119773
rect 186281 119745 186309 119773
rect 201579 119931 201607 119959
rect 201641 119931 201669 119959
rect 201579 119869 201607 119897
rect 201641 119869 201669 119897
rect 201579 119807 201607 119835
rect 201641 119807 201669 119835
rect 201579 119745 201607 119773
rect 201641 119745 201669 119773
rect 216939 119931 216967 119959
rect 217001 119931 217029 119959
rect 216939 119869 216967 119897
rect 217001 119869 217029 119897
rect 216939 119807 216967 119835
rect 217001 119807 217029 119835
rect 216939 119745 216967 119773
rect 217001 119745 217029 119773
rect 232299 119931 232327 119959
rect 232361 119931 232389 119959
rect 232299 119869 232327 119897
rect 232361 119869 232389 119897
rect 232299 119807 232327 119835
rect 232361 119807 232389 119835
rect 232299 119745 232327 119773
rect 232361 119745 232389 119773
rect 247659 119931 247687 119959
rect 247721 119931 247749 119959
rect 247659 119869 247687 119897
rect 247721 119869 247749 119897
rect 247659 119807 247687 119835
rect 247721 119807 247749 119835
rect 247659 119745 247687 119773
rect 247721 119745 247749 119773
rect 254577 119931 254605 119959
rect 254639 119931 254667 119959
rect 254701 119931 254729 119959
rect 254763 119931 254791 119959
rect 254577 119869 254605 119897
rect 254639 119869 254667 119897
rect 254701 119869 254729 119897
rect 254763 119869 254791 119897
rect 254577 119807 254605 119835
rect 254639 119807 254667 119835
rect 254701 119807 254729 119835
rect 254763 119807 254791 119835
rect 254577 119745 254605 119773
rect 254639 119745 254667 119773
rect 254701 119745 254729 119773
rect 254763 119745 254791 119773
rect 31437 113931 31465 113959
rect 31499 113931 31527 113959
rect 31561 113931 31589 113959
rect 31623 113931 31651 113959
rect 31437 113869 31465 113897
rect 31499 113869 31527 113897
rect 31561 113869 31589 113897
rect 31623 113869 31651 113897
rect 31437 113807 31465 113835
rect 31499 113807 31527 113835
rect 31561 113807 31589 113835
rect 31623 113807 31651 113835
rect 31437 113745 31465 113773
rect 31499 113745 31527 113773
rect 31561 113745 31589 113773
rect 31623 113745 31651 113773
rect 40299 113931 40327 113959
rect 40361 113931 40389 113959
rect 40299 113869 40327 113897
rect 40361 113869 40389 113897
rect 40299 113807 40327 113835
rect 40361 113807 40389 113835
rect 40299 113745 40327 113773
rect 40361 113745 40389 113773
rect 55659 113931 55687 113959
rect 55721 113931 55749 113959
rect 55659 113869 55687 113897
rect 55721 113869 55749 113897
rect 55659 113807 55687 113835
rect 55721 113807 55749 113835
rect 55659 113745 55687 113773
rect 55721 113745 55749 113773
rect 71019 113931 71047 113959
rect 71081 113931 71109 113959
rect 71019 113869 71047 113897
rect 71081 113869 71109 113897
rect 71019 113807 71047 113835
rect 71081 113807 71109 113835
rect 71019 113745 71047 113773
rect 71081 113745 71109 113773
rect 86379 113931 86407 113959
rect 86441 113931 86469 113959
rect 86379 113869 86407 113897
rect 86441 113869 86469 113897
rect 86379 113807 86407 113835
rect 86441 113807 86469 113835
rect 86379 113745 86407 113773
rect 86441 113745 86469 113773
rect 101739 113931 101767 113959
rect 101801 113931 101829 113959
rect 101739 113869 101767 113897
rect 101801 113869 101829 113897
rect 101739 113807 101767 113835
rect 101801 113807 101829 113835
rect 101739 113745 101767 113773
rect 101801 113745 101829 113773
rect 117099 113931 117127 113959
rect 117161 113931 117189 113959
rect 117099 113869 117127 113897
rect 117161 113869 117189 113897
rect 117099 113807 117127 113835
rect 117161 113807 117189 113835
rect 117099 113745 117127 113773
rect 117161 113745 117189 113773
rect 132459 113931 132487 113959
rect 132521 113931 132549 113959
rect 132459 113869 132487 113897
rect 132521 113869 132549 113897
rect 132459 113807 132487 113835
rect 132521 113807 132549 113835
rect 132459 113745 132487 113773
rect 132521 113745 132549 113773
rect 147819 113931 147847 113959
rect 147881 113931 147909 113959
rect 147819 113869 147847 113897
rect 147881 113869 147909 113897
rect 147819 113807 147847 113835
rect 147881 113807 147909 113835
rect 147819 113745 147847 113773
rect 147881 113745 147909 113773
rect 163179 113931 163207 113959
rect 163241 113931 163269 113959
rect 163179 113869 163207 113897
rect 163241 113869 163269 113897
rect 163179 113807 163207 113835
rect 163241 113807 163269 113835
rect 163179 113745 163207 113773
rect 163241 113745 163269 113773
rect 178539 113931 178567 113959
rect 178601 113931 178629 113959
rect 178539 113869 178567 113897
rect 178601 113869 178629 113897
rect 178539 113807 178567 113835
rect 178601 113807 178629 113835
rect 178539 113745 178567 113773
rect 178601 113745 178629 113773
rect 193899 113931 193927 113959
rect 193961 113931 193989 113959
rect 193899 113869 193927 113897
rect 193961 113869 193989 113897
rect 193899 113807 193927 113835
rect 193961 113807 193989 113835
rect 193899 113745 193927 113773
rect 193961 113745 193989 113773
rect 209259 113931 209287 113959
rect 209321 113931 209349 113959
rect 209259 113869 209287 113897
rect 209321 113869 209349 113897
rect 209259 113807 209287 113835
rect 209321 113807 209349 113835
rect 209259 113745 209287 113773
rect 209321 113745 209349 113773
rect 224619 113931 224647 113959
rect 224681 113931 224709 113959
rect 224619 113869 224647 113897
rect 224681 113869 224709 113897
rect 224619 113807 224647 113835
rect 224681 113807 224709 113835
rect 224619 113745 224647 113773
rect 224681 113745 224709 113773
rect 239979 113931 240007 113959
rect 240041 113931 240069 113959
rect 239979 113869 240007 113897
rect 240041 113869 240069 113897
rect 239979 113807 240007 113835
rect 240041 113807 240069 113835
rect 239979 113745 240007 113773
rect 240041 113745 240069 113773
rect 32619 110931 32647 110959
rect 32681 110931 32709 110959
rect 32619 110869 32647 110897
rect 32681 110869 32709 110897
rect 32619 110807 32647 110835
rect 32681 110807 32709 110835
rect 32619 110745 32647 110773
rect 32681 110745 32709 110773
rect 47979 110931 48007 110959
rect 48041 110931 48069 110959
rect 47979 110869 48007 110897
rect 48041 110869 48069 110897
rect 47979 110807 48007 110835
rect 48041 110807 48069 110835
rect 47979 110745 48007 110773
rect 48041 110745 48069 110773
rect 63339 110931 63367 110959
rect 63401 110931 63429 110959
rect 63339 110869 63367 110897
rect 63401 110869 63429 110897
rect 63339 110807 63367 110835
rect 63401 110807 63429 110835
rect 63339 110745 63367 110773
rect 63401 110745 63429 110773
rect 78699 110931 78727 110959
rect 78761 110931 78789 110959
rect 78699 110869 78727 110897
rect 78761 110869 78789 110897
rect 78699 110807 78727 110835
rect 78761 110807 78789 110835
rect 78699 110745 78727 110773
rect 78761 110745 78789 110773
rect 94059 110931 94087 110959
rect 94121 110931 94149 110959
rect 94059 110869 94087 110897
rect 94121 110869 94149 110897
rect 94059 110807 94087 110835
rect 94121 110807 94149 110835
rect 94059 110745 94087 110773
rect 94121 110745 94149 110773
rect 109419 110931 109447 110959
rect 109481 110931 109509 110959
rect 109419 110869 109447 110897
rect 109481 110869 109509 110897
rect 109419 110807 109447 110835
rect 109481 110807 109509 110835
rect 109419 110745 109447 110773
rect 109481 110745 109509 110773
rect 124779 110931 124807 110959
rect 124841 110931 124869 110959
rect 124779 110869 124807 110897
rect 124841 110869 124869 110897
rect 124779 110807 124807 110835
rect 124841 110807 124869 110835
rect 124779 110745 124807 110773
rect 124841 110745 124869 110773
rect 140139 110931 140167 110959
rect 140201 110931 140229 110959
rect 140139 110869 140167 110897
rect 140201 110869 140229 110897
rect 140139 110807 140167 110835
rect 140201 110807 140229 110835
rect 140139 110745 140167 110773
rect 140201 110745 140229 110773
rect 155499 110931 155527 110959
rect 155561 110931 155589 110959
rect 155499 110869 155527 110897
rect 155561 110869 155589 110897
rect 155499 110807 155527 110835
rect 155561 110807 155589 110835
rect 155499 110745 155527 110773
rect 155561 110745 155589 110773
rect 170859 110931 170887 110959
rect 170921 110931 170949 110959
rect 170859 110869 170887 110897
rect 170921 110869 170949 110897
rect 170859 110807 170887 110835
rect 170921 110807 170949 110835
rect 170859 110745 170887 110773
rect 170921 110745 170949 110773
rect 186219 110931 186247 110959
rect 186281 110931 186309 110959
rect 186219 110869 186247 110897
rect 186281 110869 186309 110897
rect 186219 110807 186247 110835
rect 186281 110807 186309 110835
rect 186219 110745 186247 110773
rect 186281 110745 186309 110773
rect 201579 110931 201607 110959
rect 201641 110931 201669 110959
rect 201579 110869 201607 110897
rect 201641 110869 201669 110897
rect 201579 110807 201607 110835
rect 201641 110807 201669 110835
rect 201579 110745 201607 110773
rect 201641 110745 201669 110773
rect 216939 110931 216967 110959
rect 217001 110931 217029 110959
rect 216939 110869 216967 110897
rect 217001 110869 217029 110897
rect 216939 110807 216967 110835
rect 217001 110807 217029 110835
rect 216939 110745 216967 110773
rect 217001 110745 217029 110773
rect 232299 110931 232327 110959
rect 232361 110931 232389 110959
rect 232299 110869 232327 110897
rect 232361 110869 232389 110897
rect 232299 110807 232327 110835
rect 232361 110807 232389 110835
rect 232299 110745 232327 110773
rect 232361 110745 232389 110773
rect 247659 110931 247687 110959
rect 247721 110931 247749 110959
rect 247659 110869 247687 110897
rect 247721 110869 247749 110897
rect 247659 110807 247687 110835
rect 247721 110807 247749 110835
rect 247659 110745 247687 110773
rect 247721 110745 247749 110773
rect 254577 110931 254605 110959
rect 254639 110931 254667 110959
rect 254701 110931 254729 110959
rect 254763 110931 254791 110959
rect 254577 110869 254605 110897
rect 254639 110869 254667 110897
rect 254701 110869 254729 110897
rect 254763 110869 254791 110897
rect 254577 110807 254605 110835
rect 254639 110807 254667 110835
rect 254701 110807 254729 110835
rect 254763 110807 254791 110835
rect 254577 110745 254605 110773
rect 254639 110745 254667 110773
rect 254701 110745 254729 110773
rect 254763 110745 254791 110773
rect 31437 104931 31465 104959
rect 31499 104931 31527 104959
rect 31561 104931 31589 104959
rect 31623 104931 31651 104959
rect 31437 104869 31465 104897
rect 31499 104869 31527 104897
rect 31561 104869 31589 104897
rect 31623 104869 31651 104897
rect 31437 104807 31465 104835
rect 31499 104807 31527 104835
rect 31561 104807 31589 104835
rect 31623 104807 31651 104835
rect 31437 104745 31465 104773
rect 31499 104745 31527 104773
rect 31561 104745 31589 104773
rect 31623 104745 31651 104773
rect 40299 104931 40327 104959
rect 40361 104931 40389 104959
rect 40299 104869 40327 104897
rect 40361 104869 40389 104897
rect 40299 104807 40327 104835
rect 40361 104807 40389 104835
rect 40299 104745 40327 104773
rect 40361 104745 40389 104773
rect 55659 104931 55687 104959
rect 55721 104931 55749 104959
rect 55659 104869 55687 104897
rect 55721 104869 55749 104897
rect 55659 104807 55687 104835
rect 55721 104807 55749 104835
rect 55659 104745 55687 104773
rect 55721 104745 55749 104773
rect 71019 104931 71047 104959
rect 71081 104931 71109 104959
rect 71019 104869 71047 104897
rect 71081 104869 71109 104897
rect 71019 104807 71047 104835
rect 71081 104807 71109 104835
rect 71019 104745 71047 104773
rect 71081 104745 71109 104773
rect 86379 104931 86407 104959
rect 86441 104931 86469 104959
rect 86379 104869 86407 104897
rect 86441 104869 86469 104897
rect 86379 104807 86407 104835
rect 86441 104807 86469 104835
rect 86379 104745 86407 104773
rect 86441 104745 86469 104773
rect 101739 104931 101767 104959
rect 101801 104931 101829 104959
rect 101739 104869 101767 104897
rect 101801 104869 101829 104897
rect 101739 104807 101767 104835
rect 101801 104807 101829 104835
rect 101739 104745 101767 104773
rect 101801 104745 101829 104773
rect 117099 104931 117127 104959
rect 117161 104931 117189 104959
rect 117099 104869 117127 104897
rect 117161 104869 117189 104897
rect 117099 104807 117127 104835
rect 117161 104807 117189 104835
rect 117099 104745 117127 104773
rect 117161 104745 117189 104773
rect 132459 104931 132487 104959
rect 132521 104931 132549 104959
rect 132459 104869 132487 104897
rect 132521 104869 132549 104897
rect 132459 104807 132487 104835
rect 132521 104807 132549 104835
rect 132459 104745 132487 104773
rect 132521 104745 132549 104773
rect 147819 104931 147847 104959
rect 147881 104931 147909 104959
rect 147819 104869 147847 104897
rect 147881 104869 147909 104897
rect 147819 104807 147847 104835
rect 147881 104807 147909 104835
rect 147819 104745 147847 104773
rect 147881 104745 147909 104773
rect 163179 104931 163207 104959
rect 163241 104931 163269 104959
rect 163179 104869 163207 104897
rect 163241 104869 163269 104897
rect 163179 104807 163207 104835
rect 163241 104807 163269 104835
rect 163179 104745 163207 104773
rect 163241 104745 163269 104773
rect 178539 104931 178567 104959
rect 178601 104931 178629 104959
rect 178539 104869 178567 104897
rect 178601 104869 178629 104897
rect 178539 104807 178567 104835
rect 178601 104807 178629 104835
rect 178539 104745 178567 104773
rect 178601 104745 178629 104773
rect 193899 104931 193927 104959
rect 193961 104931 193989 104959
rect 193899 104869 193927 104897
rect 193961 104869 193989 104897
rect 193899 104807 193927 104835
rect 193961 104807 193989 104835
rect 193899 104745 193927 104773
rect 193961 104745 193989 104773
rect 209259 104931 209287 104959
rect 209321 104931 209349 104959
rect 209259 104869 209287 104897
rect 209321 104869 209349 104897
rect 209259 104807 209287 104835
rect 209321 104807 209349 104835
rect 209259 104745 209287 104773
rect 209321 104745 209349 104773
rect 224619 104931 224647 104959
rect 224681 104931 224709 104959
rect 224619 104869 224647 104897
rect 224681 104869 224709 104897
rect 224619 104807 224647 104835
rect 224681 104807 224709 104835
rect 224619 104745 224647 104773
rect 224681 104745 224709 104773
rect 239979 104931 240007 104959
rect 240041 104931 240069 104959
rect 239979 104869 240007 104897
rect 240041 104869 240069 104897
rect 239979 104807 240007 104835
rect 240041 104807 240069 104835
rect 239979 104745 240007 104773
rect 240041 104745 240069 104773
rect 32619 101931 32647 101959
rect 32681 101931 32709 101959
rect 32619 101869 32647 101897
rect 32681 101869 32709 101897
rect 32619 101807 32647 101835
rect 32681 101807 32709 101835
rect 32619 101745 32647 101773
rect 32681 101745 32709 101773
rect 47979 101931 48007 101959
rect 48041 101931 48069 101959
rect 47979 101869 48007 101897
rect 48041 101869 48069 101897
rect 47979 101807 48007 101835
rect 48041 101807 48069 101835
rect 47979 101745 48007 101773
rect 48041 101745 48069 101773
rect 63339 101931 63367 101959
rect 63401 101931 63429 101959
rect 63339 101869 63367 101897
rect 63401 101869 63429 101897
rect 63339 101807 63367 101835
rect 63401 101807 63429 101835
rect 63339 101745 63367 101773
rect 63401 101745 63429 101773
rect 78699 101931 78727 101959
rect 78761 101931 78789 101959
rect 78699 101869 78727 101897
rect 78761 101869 78789 101897
rect 78699 101807 78727 101835
rect 78761 101807 78789 101835
rect 78699 101745 78727 101773
rect 78761 101745 78789 101773
rect 94059 101931 94087 101959
rect 94121 101931 94149 101959
rect 94059 101869 94087 101897
rect 94121 101869 94149 101897
rect 94059 101807 94087 101835
rect 94121 101807 94149 101835
rect 94059 101745 94087 101773
rect 94121 101745 94149 101773
rect 109419 101931 109447 101959
rect 109481 101931 109509 101959
rect 109419 101869 109447 101897
rect 109481 101869 109509 101897
rect 109419 101807 109447 101835
rect 109481 101807 109509 101835
rect 109419 101745 109447 101773
rect 109481 101745 109509 101773
rect 124779 101931 124807 101959
rect 124841 101931 124869 101959
rect 124779 101869 124807 101897
rect 124841 101869 124869 101897
rect 124779 101807 124807 101835
rect 124841 101807 124869 101835
rect 124779 101745 124807 101773
rect 124841 101745 124869 101773
rect 140139 101931 140167 101959
rect 140201 101931 140229 101959
rect 140139 101869 140167 101897
rect 140201 101869 140229 101897
rect 140139 101807 140167 101835
rect 140201 101807 140229 101835
rect 140139 101745 140167 101773
rect 140201 101745 140229 101773
rect 155499 101931 155527 101959
rect 155561 101931 155589 101959
rect 155499 101869 155527 101897
rect 155561 101869 155589 101897
rect 155499 101807 155527 101835
rect 155561 101807 155589 101835
rect 155499 101745 155527 101773
rect 155561 101745 155589 101773
rect 170859 101931 170887 101959
rect 170921 101931 170949 101959
rect 170859 101869 170887 101897
rect 170921 101869 170949 101897
rect 170859 101807 170887 101835
rect 170921 101807 170949 101835
rect 170859 101745 170887 101773
rect 170921 101745 170949 101773
rect 186219 101931 186247 101959
rect 186281 101931 186309 101959
rect 186219 101869 186247 101897
rect 186281 101869 186309 101897
rect 186219 101807 186247 101835
rect 186281 101807 186309 101835
rect 186219 101745 186247 101773
rect 186281 101745 186309 101773
rect 201579 101931 201607 101959
rect 201641 101931 201669 101959
rect 201579 101869 201607 101897
rect 201641 101869 201669 101897
rect 201579 101807 201607 101835
rect 201641 101807 201669 101835
rect 201579 101745 201607 101773
rect 201641 101745 201669 101773
rect 216939 101931 216967 101959
rect 217001 101931 217029 101959
rect 216939 101869 216967 101897
rect 217001 101869 217029 101897
rect 216939 101807 216967 101835
rect 217001 101807 217029 101835
rect 216939 101745 216967 101773
rect 217001 101745 217029 101773
rect 232299 101931 232327 101959
rect 232361 101931 232389 101959
rect 232299 101869 232327 101897
rect 232361 101869 232389 101897
rect 232299 101807 232327 101835
rect 232361 101807 232389 101835
rect 232299 101745 232327 101773
rect 232361 101745 232389 101773
rect 247659 101931 247687 101959
rect 247721 101931 247749 101959
rect 247659 101869 247687 101897
rect 247721 101869 247749 101897
rect 247659 101807 247687 101835
rect 247721 101807 247749 101835
rect 247659 101745 247687 101773
rect 247721 101745 247749 101773
rect 254577 101931 254605 101959
rect 254639 101931 254667 101959
rect 254701 101931 254729 101959
rect 254763 101931 254791 101959
rect 254577 101869 254605 101897
rect 254639 101869 254667 101897
rect 254701 101869 254729 101897
rect 254763 101869 254791 101897
rect 254577 101807 254605 101835
rect 254639 101807 254667 101835
rect 254701 101807 254729 101835
rect 254763 101807 254791 101835
rect 254577 101745 254605 101773
rect 254639 101745 254667 101773
rect 254701 101745 254729 101773
rect 254763 101745 254791 101773
rect 31437 95931 31465 95959
rect 31499 95931 31527 95959
rect 31561 95931 31589 95959
rect 31623 95931 31651 95959
rect 31437 95869 31465 95897
rect 31499 95869 31527 95897
rect 31561 95869 31589 95897
rect 31623 95869 31651 95897
rect 31437 95807 31465 95835
rect 31499 95807 31527 95835
rect 31561 95807 31589 95835
rect 31623 95807 31651 95835
rect 31437 95745 31465 95773
rect 31499 95745 31527 95773
rect 31561 95745 31589 95773
rect 31623 95745 31651 95773
rect 40299 95931 40327 95959
rect 40361 95931 40389 95959
rect 40299 95869 40327 95897
rect 40361 95869 40389 95897
rect 40299 95807 40327 95835
rect 40361 95807 40389 95835
rect 40299 95745 40327 95773
rect 40361 95745 40389 95773
rect 55659 95931 55687 95959
rect 55721 95931 55749 95959
rect 55659 95869 55687 95897
rect 55721 95869 55749 95897
rect 55659 95807 55687 95835
rect 55721 95807 55749 95835
rect 55659 95745 55687 95773
rect 55721 95745 55749 95773
rect 71019 95931 71047 95959
rect 71081 95931 71109 95959
rect 71019 95869 71047 95897
rect 71081 95869 71109 95897
rect 71019 95807 71047 95835
rect 71081 95807 71109 95835
rect 71019 95745 71047 95773
rect 71081 95745 71109 95773
rect 86379 95931 86407 95959
rect 86441 95931 86469 95959
rect 86379 95869 86407 95897
rect 86441 95869 86469 95897
rect 86379 95807 86407 95835
rect 86441 95807 86469 95835
rect 86379 95745 86407 95773
rect 86441 95745 86469 95773
rect 101739 95931 101767 95959
rect 101801 95931 101829 95959
rect 101739 95869 101767 95897
rect 101801 95869 101829 95897
rect 101739 95807 101767 95835
rect 101801 95807 101829 95835
rect 101739 95745 101767 95773
rect 101801 95745 101829 95773
rect 117099 95931 117127 95959
rect 117161 95931 117189 95959
rect 117099 95869 117127 95897
rect 117161 95869 117189 95897
rect 117099 95807 117127 95835
rect 117161 95807 117189 95835
rect 117099 95745 117127 95773
rect 117161 95745 117189 95773
rect 132459 95931 132487 95959
rect 132521 95931 132549 95959
rect 132459 95869 132487 95897
rect 132521 95869 132549 95897
rect 132459 95807 132487 95835
rect 132521 95807 132549 95835
rect 132459 95745 132487 95773
rect 132521 95745 132549 95773
rect 147819 95931 147847 95959
rect 147881 95931 147909 95959
rect 147819 95869 147847 95897
rect 147881 95869 147909 95897
rect 147819 95807 147847 95835
rect 147881 95807 147909 95835
rect 147819 95745 147847 95773
rect 147881 95745 147909 95773
rect 163179 95931 163207 95959
rect 163241 95931 163269 95959
rect 163179 95869 163207 95897
rect 163241 95869 163269 95897
rect 163179 95807 163207 95835
rect 163241 95807 163269 95835
rect 163179 95745 163207 95773
rect 163241 95745 163269 95773
rect 178539 95931 178567 95959
rect 178601 95931 178629 95959
rect 178539 95869 178567 95897
rect 178601 95869 178629 95897
rect 178539 95807 178567 95835
rect 178601 95807 178629 95835
rect 178539 95745 178567 95773
rect 178601 95745 178629 95773
rect 193899 95931 193927 95959
rect 193961 95931 193989 95959
rect 193899 95869 193927 95897
rect 193961 95869 193989 95897
rect 193899 95807 193927 95835
rect 193961 95807 193989 95835
rect 193899 95745 193927 95773
rect 193961 95745 193989 95773
rect 209259 95931 209287 95959
rect 209321 95931 209349 95959
rect 209259 95869 209287 95897
rect 209321 95869 209349 95897
rect 209259 95807 209287 95835
rect 209321 95807 209349 95835
rect 209259 95745 209287 95773
rect 209321 95745 209349 95773
rect 224619 95931 224647 95959
rect 224681 95931 224709 95959
rect 224619 95869 224647 95897
rect 224681 95869 224709 95897
rect 224619 95807 224647 95835
rect 224681 95807 224709 95835
rect 224619 95745 224647 95773
rect 224681 95745 224709 95773
rect 239979 95931 240007 95959
rect 240041 95931 240069 95959
rect 239979 95869 240007 95897
rect 240041 95869 240069 95897
rect 239979 95807 240007 95835
rect 240041 95807 240069 95835
rect 239979 95745 240007 95773
rect 240041 95745 240069 95773
rect 32619 92931 32647 92959
rect 32681 92931 32709 92959
rect 32619 92869 32647 92897
rect 32681 92869 32709 92897
rect 32619 92807 32647 92835
rect 32681 92807 32709 92835
rect 32619 92745 32647 92773
rect 32681 92745 32709 92773
rect 47979 92931 48007 92959
rect 48041 92931 48069 92959
rect 47979 92869 48007 92897
rect 48041 92869 48069 92897
rect 47979 92807 48007 92835
rect 48041 92807 48069 92835
rect 47979 92745 48007 92773
rect 48041 92745 48069 92773
rect 63339 92931 63367 92959
rect 63401 92931 63429 92959
rect 63339 92869 63367 92897
rect 63401 92869 63429 92897
rect 63339 92807 63367 92835
rect 63401 92807 63429 92835
rect 63339 92745 63367 92773
rect 63401 92745 63429 92773
rect 78699 92931 78727 92959
rect 78761 92931 78789 92959
rect 78699 92869 78727 92897
rect 78761 92869 78789 92897
rect 78699 92807 78727 92835
rect 78761 92807 78789 92835
rect 78699 92745 78727 92773
rect 78761 92745 78789 92773
rect 94059 92931 94087 92959
rect 94121 92931 94149 92959
rect 94059 92869 94087 92897
rect 94121 92869 94149 92897
rect 94059 92807 94087 92835
rect 94121 92807 94149 92835
rect 94059 92745 94087 92773
rect 94121 92745 94149 92773
rect 109419 92931 109447 92959
rect 109481 92931 109509 92959
rect 109419 92869 109447 92897
rect 109481 92869 109509 92897
rect 109419 92807 109447 92835
rect 109481 92807 109509 92835
rect 109419 92745 109447 92773
rect 109481 92745 109509 92773
rect 124779 92931 124807 92959
rect 124841 92931 124869 92959
rect 124779 92869 124807 92897
rect 124841 92869 124869 92897
rect 124779 92807 124807 92835
rect 124841 92807 124869 92835
rect 124779 92745 124807 92773
rect 124841 92745 124869 92773
rect 140139 92931 140167 92959
rect 140201 92931 140229 92959
rect 140139 92869 140167 92897
rect 140201 92869 140229 92897
rect 140139 92807 140167 92835
rect 140201 92807 140229 92835
rect 140139 92745 140167 92773
rect 140201 92745 140229 92773
rect 155499 92931 155527 92959
rect 155561 92931 155589 92959
rect 155499 92869 155527 92897
rect 155561 92869 155589 92897
rect 155499 92807 155527 92835
rect 155561 92807 155589 92835
rect 155499 92745 155527 92773
rect 155561 92745 155589 92773
rect 170859 92931 170887 92959
rect 170921 92931 170949 92959
rect 170859 92869 170887 92897
rect 170921 92869 170949 92897
rect 170859 92807 170887 92835
rect 170921 92807 170949 92835
rect 170859 92745 170887 92773
rect 170921 92745 170949 92773
rect 186219 92931 186247 92959
rect 186281 92931 186309 92959
rect 186219 92869 186247 92897
rect 186281 92869 186309 92897
rect 186219 92807 186247 92835
rect 186281 92807 186309 92835
rect 186219 92745 186247 92773
rect 186281 92745 186309 92773
rect 201579 92931 201607 92959
rect 201641 92931 201669 92959
rect 201579 92869 201607 92897
rect 201641 92869 201669 92897
rect 201579 92807 201607 92835
rect 201641 92807 201669 92835
rect 201579 92745 201607 92773
rect 201641 92745 201669 92773
rect 216939 92931 216967 92959
rect 217001 92931 217029 92959
rect 216939 92869 216967 92897
rect 217001 92869 217029 92897
rect 216939 92807 216967 92835
rect 217001 92807 217029 92835
rect 216939 92745 216967 92773
rect 217001 92745 217029 92773
rect 232299 92931 232327 92959
rect 232361 92931 232389 92959
rect 232299 92869 232327 92897
rect 232361 92869 232389 92897
rect 232299 92807 232327 92835
rect 232361 92807 232389 92835
rect 232299 92745 232327 92773
rect 232361 92745 232389 92773
rect 247659 92931 247687 92959
rect 247721 92931 247749 92959
rect 247659 92869 247687 92897
rect 247721 92869 247749 92897
rect 247659 92807 247687 92835
rect 247721 92807 247749 92835
rect 247659 92745 247687 92773
rect 247721 92745 247749 92773
rect 254577 92931 254605 92959
rect 254639 92931 254667 92959
rect 254701 92931 254729 92959
rect 254763 92931 254791 92959
rect 254577 92869 254605 92897
rect 254639 92869 254667 92897
rect 254701 92869 254729 92897
rect 254763 92869 254791 92897
rect 254577 92807 254605 92835
rect 254639 92807 254667 92835
rect 254701 92807 254729 92835
rect 254763 92807 254791 92835
rect 254577 92745 254605 92773
rect 254639 92745 254667 92773
rect 254701 92745 254729 92773
rect 254763 92745 254791 92773
rect 31437 86931 31465 86959
rect 31499 86931 31527 86959
rect 31561 86931 31589 86959
rect 31623 86931 31651 86959
rect 31437 86869 31465 86897
rect 31499 86869 31527 86897
rect 31561 86869 31589 86897
rect 31623 86869 31651 86897
rect 31437 86807 31465 86835
rect 31499 86807 31527 86835
rect 31561 86807 31589 86835
rect 31623 86807 31651 86835
rect 31437 86745 31465 86773
rect 31499 86745 31527 86773
rect 31561 86745 31589 86773
rect 31623 86745 31651 86773
rect 40299 86931 40327 86959
rect 40361 86931 40389 86959
rect 40299 86869 40327 86897
rect 40361 86869 40389 86897
rect 40299 86807 40327 86835
rect 40361 86807 40389 86835
rect 40299 86745 40327 86773
rect 40361 86745 40389 86773
rect 55659 86931 55687 86959
rect 55721 86931 55749 86959
rect 55659 86869 55687 86897
rect 55721 86869 55749 86897
rect 55659 86807 55687 86835
rect 55721 86807 55749 86835
rect 55659 86745 55687 86773
rect 55721 86745 55749 86773
rect 71019 86931 71047 86959
rect 71081 86931 71109 86959
rect 71019 86869 71047 86897
rect 71081 86869 71109 86897
rect 71019 86807 71047 86835
rect 71081 86807 71109 86835
rect 71019 86745 71047 86773
rect 71081 86745 71109 86773
rect 86379 86931 86407 86959
rect 86441 86931 86469 86959
rect 86379 86869 86407 86897
rect 86441 86869 86469 86897
rect 86379 86807 86407 86835
rect 86441 86807 86469 86835
rect 86379 86745 86407 86773
rect 86441 86745 86469 86773
rect 101739 86931 101767 86959
rect 101801 86931 101829 86959
rect 101739 86869 101767 86897
rect 101801 86869 101829 86897
rect 101739 86807 101767 86835
rect 101801 86807 101829 86835
rect 101739 86745 101767 86773
rect 101801 86745 101829 86773
rect 117099 86931 117127 86959
rect 117161 86931 117189 86959
rect 117099 86869 117127 86897
rect 117161 86869 117189 86897
rect 117099 86807 117127 86835
rect 117161 86807 117189 86835
rect 117099 86745 117127 86773
rect 117161 86745 117189 86773
rect 132459 86931 132487 86959
rect 132521 86931 132549 86959
rect 132459 86869 132487 86897
rect 132521 86869 132549 86897
rect 132459 86807 132487 86835
rect 132521 86807 132549 86835
rect 132459 86745 132487 86773
rect 132521 86745 132549 86773
rect 147819 86931 147847 86959
rect 147881 86931 147909 86959
rect 147819 86869 147847 86897
rect 147881 86869 147909 86897
rect 147819 86807 147847 86835
rect 147881 86807 147909 86835
rect 147819 86745 147847 86773
rect 147881 86745 147909 86773
rect 163179 86931 163207 86959
rect 163241 86931 163269 86959
rect 163179 86869 163207 86897
rect 163241 86869 163269 86897
rect 163179 86807 163207 86835
rect 163241 86807 163269 86835
rect 163179 86745 163207 86773
rect 163241 86745 163269 86773
rect 178539 86931 178567 86959
rect 178601 86931 178629 86959
rect 178539 86869 178567 86897
rect 178601 86869 178629 86897
rect 178539 86807 178567 86835
rect 178601 86807 178629 86835
rect 178539 86745 178567 86773
rect 178601 86745 178629 86773
rect 193899 86931 193927 86959
rect 193961 86931 193989 86959
rect 193899 86869 193927 86897
rect 193961 86869 193989 86897
rect 193899 86807 193927 86835
rect 193961 86807 193989 86835
rect 193899 86745 193927 86773
rect 193961 86745 193989 86773
rect 209259 86931 209287 86959
rect 209321 86931 209349 86959
rect 209259 86869 209287 86897
rect 209321 86869 209349 86897
rect 209259 86807 209287 86835
rect 209321 86807 209349 86835
rect 209259 86745 209287 86773
rect 209321 86745 209349 86773
rect 224619 86931 224647 86959
rect 224681 86931 224709 86959
rect 224619 86869 224647 86897
rect 224681 86869 224709 86897
rect 224619 86807 224647 86835
rect 224681 86807 224709 86835
rect 224619 86745 224647 86773
rect 224681 86745 224709 86773
rect 239979 86931 240007 86959
rect 240041 86931 240069 86959
rect 239979 86869 240007 86897
rect 240041 86869 240069 86897
rect 239979 86807 240007 86835
rect 240041 86807 240069 86835
rect 239979 86745 240007 86773
rect 240041 86745 240069 86773
rect 32619 83931 32647 83959
rect 32681 83931 32709 83959
rect 32619 83869 32647 83897
rect 32681 83869 32709 83897
rect 32619 83807 32647 83835
rect 32681 83807 32709 83835
rect 32619 83745 32647 83773
rect 32681 83745 32709 83773
rect 47979 83931 48007 83959
rect 48041 83931 48069 83959
rect 47979 83869 48007 83897
rect 48041 83869 48069 83897
rect 47979 83807 48007 83835
rect 48041 83807 48069 83835
rect 47979 83745 48007 83773
rect 48041 83745 48069 83773
rect 63339 83931 63367 83959
rect 63401 83931 63429 83959
rect 63339 83869 63367 83897
rect 63401 83869 63429 83897
rect 63339 83807 63367 83835
rect 63401 83807 63429 83835
rect 63339 83745 63367 83773
rect 63401 83745 63429 83773
rect 78699 83931 78727 83959
rect 78761 83931 78789 83959
rect 78699 83869 78727 83897
rect 78761 83869 78789 83897
rect 78699 83807 78727 83835
rect 78761 83807 78789 83835
rect 78699 83745 78727 83773
rect 78761 83745 78789 83773
rect 94059 83931 94087 83959
rect 94121 83931 94149 83959
rect 94059 83869 94087 83897
rect 94121 83869 94149 83897
rect 94059 83807 94087 83835
rect 94121 83807 94149 83835
rect 94059 83745 94087 83773
rect 94121 83745 94149 83773
rect 109419 83931 109447 83959
rect 109481 83931 109509 83959
rect 109419 83869 109447 83897
rect 109481 83869 109509 83897
rect 109419 83807 109447 83835
rect 109481 83807 109509 83835
rect 109419 83745 109447 83773
rect 109481 83745 109509 83773
rect 124779 83931 124807 83959
rect 124841 83931 124869 83959
rect 124779 83869 124807 83897
rect 124841 83869 124869 83897
rect 124779 83807 124807 83835
rect 124841 83807 124869 83835
rect 124779 83745 124807 83773
rect 124841 83745 124869 83773
rect 140139 83931 140167 83959
rect 140201 83931 140229 83959
rect 140139 83869 140167 83897
rect 140201 83869 140229 83897
rect 140139 83807 140167 83835
rect 140201 83807 140229 83835
rect 140139 83745 140167 83773
rect 140201 83745 140229 83773
rect 155499 83931 155527 83959
rect 155561 83931 155589 83959
rect 155499 83869 155527 83897
rect 155561 83869 155589 83897
rect 155499 83807 155527 83835
rect 155561 83807 155589 83835
rect 155499 83745 155527 83773
rect 155561 83745 155589 83773
rect 170859 83931 170887 83959
rect 170921 83931 170949 83959
rect 170859 83869 170887 83897
rect 170921 83869 170949 83897
rect 170859 83807 170887 83835
rect 170921 83807 170949 83835
rect 170859 83745 170887 83773
rect 170921 83745 170949 83773
rect 186219 83931 186247 83959
rect 186281 83931 186309 83959
rect 186219 83869 186247 83897
rect 186281 83869 186309 83897
rect 186219 83807 186247 83835
rect 186281 83807 186309 83835
rect 186219 83745 186247 83773
rect 186281 83745 186309 83773
rect 201579 83931 201607 83959
rect 201641 83931 201669 83959
rect 201579 83869 201607 83897
rect 201641 83869 201669 83897
rect 201579 83807 201607 83835
rect 201641 83807 201669 83835
rect 201579 83745 201607 83773
rect 201641 83745 201669 83773
rect 216939 83931 216967 83959
rect 217001 83931 217029 83959
rect 216939 83869 216967 83897
rect 217001 83869 217029 83897
rect 216939 83807 216967 83835
rect 217001 83807 217029 83835
rect 216939 83745 216967 83773
rect 217001 83745 217029 83773
rect 232299 83931 232327 83959
rect 232361 83931 232389 83959
rect 232299 83869 232327 83897
rect 232361 83869 232389 83897
rect 232299 83807 232327 83835
rect 232361 83807 232389 83835
rect 232299 83745 232327 83773
rect 232361 83745 232389 83773
rect 247659 83931 247687 83959
rect 247721 83931 247749 83959
rect 247659 83869 247687 83897
rect 247721 83869 247749 83897
rect 247659 83807 247687 83835
rect 247721 83807 247749 83835
rect 247659 83745 247687 83773
rect 247721 83745 247749 83773
rect 254577 83931 254605 83959
rect 254639 83931 254667 83959
rect 254701 83931 254729 83959
rect 254763 83931 254791 83959
rect 254577 83869 254605 83897
rect 254639 83869 254667 83897
rect 254701 83869 254729 83897
rect 254763 83869 254791 83897
rect 254577 83807 254605 83835
rect 254639 83807 254667 83835
rect 254701 83807 254729 83835
rect 254763 83807 254791 83835
rect 254577 83745 254605 83773
rect 254639 83745 254667 83773
rect 254701 83745 254729 83773
rect 254763 83745 254791 83773
rect 31437 77931 31465 77959
rect 31499 77931 31527 77959
rect 31561 77931 31589 77959
rect 31623 77931 31651 77959
rect 31437 77869 31465 77897
rect 31499 77869 31527 77897
rect 31561 77869 31589 77897
rect 31623 77869 31651 77897
rect 31437 77807 31465 77835
rect 31499 77807 31527 77835
rect 31561 77807 31589 77835
rect 31623 77807 31651 77835
rect 31437 77745 31465 77773
rect 31499 77745 31527 77773
rect 31561 77745 31589 77773
rect 31623 77745 31651 77773
rect 40299 77931 40327 77959
rect 40361 77931 40389 77959
rect 40299 77869 40327 77897
rect 40361 77869 40389 77897
rect 40299 77807 40327 77835
rect 40361 77807 40389 77835
rect 40299 77745 40327 77773
rect 40361 77745 40389 77773
rect 55659 77931 55687 77959
rect 55721 77931 55749 77959
rect 55659 77869 55687 77897
rect 55721 77869 55749 77897
rect 55659 77807 55687 77835
rect 55721 77807 55749 77835
rect 55659 77745 55687 77773
rect 55721 77745 55749 77773
rect 71019 77931 71047 77959
rect 71081 77931 71109 77959
rect 71019 77869 71047 77897
rect 71081 77869 71109 77897
rect 71019 77807 71047 77835
rect 71081 77807 71109 77835
rect 71019 77745 71047 77773
rect 71081 77745 71109 77773
rect 86379 77931 86407 77959
rect 86441 77931 86469 77959
rect 86379 77869 86407 77897
rect 86441 77869 86469 77897
rect 86379 77807 86407 77835
rect 86441 77807 86469 77835
rect 86379 77745 86407 77773
rect 86441 77745 86469 77773
rect 101739 77931 101767 77959
rect 101801 77931 101829 77959
rect 101739 77869 101767 77897
rect 101801 77869 101829 77897
rect 101739 77807 101767 77835
rect 101801 77807 101829 77835
rect 101739 77745 101767 77773
rect 101801 77745 101829 77773
rect 117099 77931 117127 77959
rect 117161 77931 117189 77959
rect 117099 77869 117127 77897
rect 117161 77869 117189 77897
rect 117099 77807 117127 77835
rect 117161 77807 117189 77835
rect 117099 77745 117127 77773
rect 117161 77745 117189 77773
rect 132459 77931 132487 77959
rect 132521 77931 132549 77959
rect 132459 77869 132487 77897
rect 132521 77869 132549 77897
rect 132459 77807 132487 77835
rect 132521 77807 132549 77835
rect 132459 77745 132487 77773
rect 132521 77745 132549 77773
rect 147819 77931 147847 77959
rect 147881 77931 147909 77959
rect 147819 77869 147847 77897
rect 147881 77869 147909 77897
rect 147819 77807 147847 77835
rect 147881 77807 147909 77835
rect 147819 77745 147847 77773
rect 147881 77745 147909 77773
rect 163179 77931 163207 77959
rect 163241 77931 163269 77959
rect 163179 77869 163207 77897
rect 163241 77869 163269 77897
rect 163179 77807 163207 77835
rect 163241 77807 163269 77835
rect 163179 77745 163207 77773
rect 163241 77745 163269 77773
rect 178539 77931 178567 77959
rect 178601 77931 178629 77959
rect 178539 77869 178567 77897
rect 178601 77869 178629 77897
rect 178539 77807 178567 77835
rect 178601 77807 178629 77835
rect 178539 77745 178567 77773
rect 178601 77745 178629 77773
rect 193899 77931 193927 77959
rect 193961 77931 193989 77959
rect 193899 77869 193927 77897
rect 193961 77869 193989 77897
rect 193899 77807 193927 77835
rect 193961 77807 193989 77835
rect 193899 77745 193927 77773
rect 193961 77745 193989 77773
rect 209259 77931 209287 77959
rect 209321 77931 209349 77959
rect 209259 77869 209287 77897
rect 209321 77869 209349 77897
rect 209259 77807 209287 77835
rect 209321 77807 209349 77835
rect 209259 77745 209287 77773
rect 209321 77745 209349 77773
rect 224619 77931 224647 77959
rect 224681 77931 224709 77959
rect 224619 77869 224647 77897
rect 224681 77869 224709 77897
rect 224619 77807 224647 77835
rect 224681 77807 224709 77835
rect 224619 77745 224647 77773
rect 224681 77745 224709 77773
rect 239979 77931 240007 77959
rect 240041 77931 240069 77959
rect 239979 77869 240007 77897
rect 240041 77869 240069 77897
rect 239979 77807 240007 77835
rect 240041 77807 240069 77835
rect 239979 77745 240007 77773
rect 240041 77745 240069 77773
rect 32619 74931 32647 74959
rect 32681 74931 32709 74959
rect 32619 74869 32647 74897
rect 32681 74869 32709 74897
rect 32619 74807 32647 74835
rect 32681 74807 32709 74835
rect 32619 74745 32647 74773
rect 32681 74745 32709 74773
rect 47979 74931 48007 74959
rect 48041 74931 48069 74959
rect 47979 74869 48007 74897
rect 48041 74869 48069 74897
rect 47979 74807 48007 74835
rect 48041 74807 48069 74835
rect 47979 74745 48007 74773
rect 48041 74745 48069 74773
rect 63339 74931 63367 74959
rect 63401 74931 63429 74959
rect 63339 74869 63367 74897
rect 63401 74869 63429 74897
rect 63339 74807 63367 74835
rect 63401 74807 63429 74835
rect 63339 74745 63367 74773
rect 63401 74745 63429 74773
rect 78699 74931 78727 74959
rect 78761 74931 78789 74959
rect 78699 74869 78727 74897
rect 78761 74869 78789 74897
rect 78699 74807 78727 74835
rect 78761 74807 78789 74835
rect 78699 74745 78727 74773
rect 78761 74745 78789 74773
rect 94059 74931 94087 74959
rect 94121 74931 94149 74959
rect 94059 74869 94087 74897
rect 94121 74869 94149 74897
rect 94059 74807 94087 74835
rect 94121 74807 94149 74835
rect 94059 74745 94087 74773
rect 94121 74745 94149 74773
rect 109419 74931 109447 74959
rect 109481 74931 109509 74959
rect 109419 74869 109447 74897
rect 109481 74869 109509 74897
rect 109419 74807 109447 74835
rect 109481 74807 109509 74835
rect 109419 74745 109447 74773
rect 109481 74745 109509 74773
rect 124779 74931 124807 74959
rect 124841 74931 124869 74959
rect 124779 74869 124807 74897
rect 124841 74869 124869 74897
rect 124779 74807 124807 74835
rect 124841 74807 124869 74835
rect 124779 74745 124807 74773
rect 124841 74745 124869 74773
rect 140139 74931 140167 74959
rect 140201 74931 140229 74959
rect 140139 74869 140167 74897
rect 140201 74869 140229 74897
rect 140139 74807 140167 74835
rect 140201 74807 140229 74835
rect 140139 74745 140167 74773
rect 140201 74745 140229 74773
rect 155499 74931 155527 74959
rect 155561 74931 155589 74959
rect 155499 74869 155527 74897
rect 155561 74869 155589 74897
rect 155499 74807 155527 74835
rect 155561 74807 155589 74835
rect 155499 74745 155527 74773
rect 155561 74745 155589 74773
rect 170859 74931 170887 74959
rect 170921 74931 170949 74959
rect 170859 74869 170887 74897
rect 170921 74869 170949 74897
rect 170859 74807 170887 74835
rect 170921 74807 170949 74835
rect 170859 74745 170887 74773
rect 170921 74745 170949 74773
rect 186219 74931 186247 74959
rect 186281 74931 186309 74959
rect 186219 74869 186247 74897
rect 186281 74869 186309 74897
rect 186219 74807 186247 74835
rect 186281 74807 186309 74835
rect 186219 74745 186247 74773
rect 186281 74745 186309 74773
rect 201579 74931 201607 74959
rect 201641 74931 201669 74959
rect 201579 74869 201607 74897
rect 201641 74869 201669 74897
rect 201579 74807 201607 74835
rect 201641 74807 201669 74835
rect 201579 74745 201607 74773
rect 201641 74745 201669 74773
rect 216939 74931 216967 74959
rect 217001 74931 217029 74959
rect 216939 74869 216967 74897
rect 217001 74869 217029 74897
rect 216939 74807 216967 74835
rect 217001 74807 217029 74835
rect 216939 74745 216967 74773
rect 217001 74745 217029 74773
rect 232299 74931 232327 74959
rect 232361 74931 232389 74959
rect 232299 74869 232327 74897
rect 232361 74869 232389 74897
rect 232299 74807 232327 74835
rect 232361 74807 232389 74835
rect 232299 74745 232327 74773
rect 232361 74745 232389 74773
rect 247659 74931 247687 74959
rect 247721 74931 247749 74959
rect 247659 74869 247687 74897
rect 247721 74869 247749 74897
rect 247659 74807 247687 74835
rect 247721 74807 247749 74835
rect 247659 74745 247687 74773
rect 247721 74745 247749 74773
rect 254577 74931 254605 74959
rect 254639 74931 254667 74959
rect 254701 74931 254729 74959
rect 254763 74931 254791 74959
rect 254577 74869 254605 74897
rect 254639 74869 254667 74897
rect 254701 74869 254729 74897
rect 254763 74869 254791 74897
rect 254577 74807 254605 74835
rect 254639 74807 254667 74835
rect 254701 74807 254729 74835
rect 254763 74807 254791 74835
rect 254577 74745 254605 74773
rect 254639 74745 254667 74773
rect 254701 74745 254729 74773
rect 254763 74745 254791 74773
rect 31437 68931 31465 68959
rect 31499 68931 31527 68959
rect 31561 68931 31589 68959
rect 31623 68931 31651 68959
rect 31437 68869 31465 68897
rect 31499 68869 31527 68897
rect 31561 68869 31589 68897
rect 31623 68869 31651 68897
rect 31437 68807 31465 68835
rect 31499 68807 31527 68835
rect 31561 68807 31589 68835
rect 31623 68807 31651 68835
rect 31437 68745 31465 68773
rect 31499 68745 31527 68773
rect 31561 68745 31589 68773
rect 31623 68745 31651 68773
rect 40299 68931 40327 68959
rect 40361 68931 40389 68959
rect 40299 68869 40327 68897
rect 40361 68869 40389 68897
rect 40299 68807 40327 68835
rect 40361 68807 40389 68835
rect 40299 68745 40327 68773
rect 40361 68745 40389 68773
rect 55659 68931 55687 68959
rect 55721 68931 55749 68959
rect 55659 68869 55687 68897
rect 55721 68869 55749 68897
rect 55659 68807 55687 68835
rect 55721 68807 55749 68835
rect 55659 68745 55687 68773
rect 55721 68745 55749 68773
rect 71019 68931 71047 68959
rect 71081 68931 71109 68959
rect 71019 68869 71047 68897
rect 71081 68869 71109 68897
rect 71019 68807 71047 68835
rect 71081 68807 71109 68835
rect 71019 68745 71047 68773
rect 71081 68745 71109 68773
rect 86379 68931 86407 68959
rect 86441 68931 86469 68959
rect 86379 68869 86407 68897
rect 86441 68869 86469 68897
rect 86379 68807 86407 68835
rect 86441 68807 86469 68835
rect 86379 68745 86407 68773
rect 86441 68745 86469 68773
rect 101739 68931 101767 68959
rect 101801 68931 101829 68959
rect 101739 68869 101767 68897
rect 101801 68869 101829 68897
rect 101739 68807 101767 68835
rect 101801 68807 101829 68835
rect 101739 68745 101767 68773
rect 101801 68745 101829 68773
rect 117099 68931 117127 68959
rect 117161 68931 117189 68959
rect 117099 68869 117127 68897
rect 117161 68869 117189 68897
rect 117099 68807 117127 68835
rect 117161 68807 117189 68835
rect 117099 68745 117127 68773
rect 117161 68745 117189 68773
rect 132459 68931 132487 68959
rect 132521 68931 132549 68959
rect 132459 68869 132487 68897
rect 132521 68869 132549 68897
rect 132459 68807 132487 68835
rect 132521 68807 132549 68835
rect 132459 68745 132487 68773
rect 132521 68745 132549 68773
rect 147819 68931 147847 68959
rect 147881 68931 147909 68959
rect 147819 68869 147847 68897
rect 147881 68869 147909 68897
rect 147819 68807 147847 68835
rect 147881 68807 147909 68835
rect 147819 68745 147847 68773
rect 147881 68745 147909 68773
rect 163179 68931 163207 68959
rect 163241 68931 163269 68959
rect 163179 68869 163207 68897
rect 163241 68869 163269 68897
rect 163179 68807 163207 68835
rect 163241 68807 163269 68835
rect 163179 68745 163207 68773
rect 163241 68745 163269 68773
rect 178539 68931 178567 68959
rect 178601 68931 178629 68959
rect 178539 68869 178567 68897
rect 178601 68869 178629 68897
rect 178539 68807 178567 68835
rect 178601 68807 178629 68835
rect 178539 68745 178567 68773
rect 178601 68745 178629 68773
rect 193899 68931 193927 68959
rect 193961 68931 193989 68959
rect 193899 68869 193927 68897
rect 193961 68869 193989 68897
rect 193899 68807 193927 68835
rect 193961 68807 193989 68835
rect 193899 68745 193927 68773
rect 193961 68745 193989 68773
rect 209259 68931 209287 68959
rect 209321 68931 209349 68959
rect 209259 68869 209287 68897
rect 209321 68869 209349 68897
rect 209259 68807 209287 68835
rect 209321 68807 209349 68835
rect 209259 68745 209287 68773
rect 209321 68745 209349 68773
rect 224619 68931 224647 68959
rect 224681 68931 224709 68959
rect 224619 68869 224647 68897
rect 224681 68869 224709 68897
rect 224619 68807 224647 68835
rect 224681 68807 224709 68835
rect 224619 68745 224647 68773
rect 224681 68745 224709 68773
rect 239979 68931 240007 68959
rect 240041 68931 240069 68959
rect 239979 68869 240007 68897
rect 240041 68869 240069 68897
rect 239979 68807 240007 68835
rect 240041 68807 240069 68835
rect 239979 68745 240007 68773
rect 240041 68745 240069 68773
rect 32619 65931 32647 65959
rect 32681 65931 32709 65959
rect 32619 65869 32647 65897
rect 32681 65869 32709 65897
rect 32619 65807 32647 65835
rect 32681 65807 32709 65835
rect 32619 65745 32647 65773
rect 32681 65745 32709 65773
rect 47979 65931 48007 65959
rect 48041 65931 48069 65959
rect 47979 65869 48007 65897
rect 48041 65869 48069 65897
rect 47979 65807 48007 65835
rect 48041 65807 48069 65835
rect 47979 65745 48007 65773
rect 48041 65745 48069 65773
rect 63339 65931 63367 65959
rect 63401 65931 63429 65959
rect 63339 65869 63367 65897
rect 63401 65869 63429 65897
rect 63339 65807 63367 65835
rect 63401 65807 63429 65835
rect 63339 65745 63367 65773
rect 63401 65745 63429 65773
rect 78699 65931 78727 65959
rect 78761 65931 78789 65959
rect 78699 65869 78727 65897
rect 78761 65869 78789 65897
rect 78699 65807 78727 65835
rect 78761 65807 78789 65835
rect 78699 65745 78727 65773
rect 78761 65745 78789 65773
rect 94059 65931 94087 65959
rect 94121 65931 94149 65959
rect 94059 65869 94087 65897
rect 94121 65869 94149 65897
rect 94059 65807 94087 65835
rect 94121 65807 94149 65835
rect 94059 65745 94087 65773
rect 94121 65745 94149 65773
rect 109419 65931 109447 65959
rect 109481 65931 109509 65959
rect 109419 65869 109447 65897
rect 109481 65869 109509 65897
rect 109419 65807 109447 65835
rect 109481 65807 109509 65835
rect 109419 65745 109447 65773
rect 109481 65745 109509 65773
rect 124779 65931 124807 65959
rect 124841 65931 124869 65959
rect 124779 65869 124807 65897
rect 124841 65869 124869 65897
rect 124779 65807 124807 65835
rect 124841 65807 124869 65835
rect 124779 65745 124807 65773
rect 124841 65745 124869 65773
rect 140139 65931 140167 65959
rect 140201 65931 140229 65959
rect 140139 65869 140167 65897
rect 140201 65869 140229 65897
rect 140139 65807 140167 65835
rect 140201 65807 140229 65835
rect 140139 65745 140167 65773
rect 140201 65745 140229 65773
rect 155499 65931 155527 65959
rect 155561 65931 155589 65959
rect 155499 65869 155527 65897
rect 155561 65869 155589 65897
rect 155499 65807 155527 65835
rect 155561 65807 155589 65835
rect 155499 65745 155527 65773
rect 155561 65745 155589 65773
rect 170859 65931 170887 65959
rect 170921 65931 170949 65959
rect 170859 65869 170887 65897
rect 170921 65869 170949 65897
rect 170859 65807 170887 65835
rect 170921 65807 170949 65835
rect 170859 65745 170887 65773
rect 170921 65745 170949 65773
rect 186219 65931 186247 65959
rect 186281 65931 186309 65959
rect 186219 65869 186247 65897
rect 186281 65869 186309 65897
rect 186219 65807 186247 65835
rect 186281 65807 186309 65835
rect 186219 65745 186247 65773
rect 186281 65745 186309 65773
rect 201579 65931 201607 65959
rect 201641 65931 201669 65959
rect 201579 65869 201607 65897
rect 201641 65869 201669 65897
rect 201579 65807 201607 65835
rect 201641 65807 201669 65835
rect 201579 65745 201607 65773
rect 201641 65745 201669 65773
rect 216939 65931 216967 65959
rect 217001 65931 217029 65959
rect 216939 65869 216967 65897
rect 217001 65869 217029 65897
rect 216939 65807 216967 65835
rect 217001 65807 217029 65835
rect 216939 65745 216967 65773
rect 217001 65745 217029 65773
rect 232299 65931 232327 65959
rect 232361 65931 232389 65959
rect 232299 65869 232327 65897
rect 232361 65869 232389 65897
rect 232299 65807 232327 65835
rect 232361 65807 232389 65835
rect 232299 65745 232327 65773
rect 232361 65745 232389 65773
rect 247659 65931 247687 65959
rect 247721 65931 247749 65959
rect 247659 65869 247687 65897
rect 247721 65869 247749 65897
rect 247659 65807 247687 65835
rect 247721 65807 247749 65835
rect 247659 65745 247687 65773
rect 247721 65745 247749 65773
rect 254577 65931 254605 65959
rect 254639 65931 254667 65959
rect 254701 65931 254729 65959
rect 254763 65931 254791 65959
rect 254577 65869 254605 65897
rect 254639 65869 254667 65897
rect 254701 65869 254729 65897
rect 254763 65869 254791 65897
rect 254577 65807 254605 65835
rect 254639 65807 254667 65835
rect 254701 65807 254729 65835
rect 254763 65807 254791 65835
rect 254577 65745 254605 65773
rect 254639 65745 254667 65773
rect 254701 65745 254729 65773
rect 254763 65745 254791 65773
rect 31437 59931 31465 59959
rect 31499 59931 31527 59959
rect 31561 59931 31589 59959
rect 31623 59931 31651 59959
rect 31437 59869 31465 59897
rect 31499 59869 31527 59897
rect 31561 59869 31589 59897
rect 31623 59869 31651 59897
rect 31437 59807 31465 59835
rect 31499 59807 31527 59835
rect 31561 59807 31589 59835
rect 31623 59807 31651 59835
rect 31437 59745 31465 59773
rect 31499 59745 31527 59773
rect 31561 59745 31589 59773
rect 31623 59745 31651 59773
rect 40299 59931 40327 59959
rect 40361 59931 40389 59959
rect 40299 59869 40327 59897
rect 40361 59869 40389 59897
rect 40299 59807 40327 59835
rect 40361 59807 40389 59835
rect 40299 59745 40327 59773
rect 40361 59745 40389 59773
rect 55659 59931 55687 59959
rect 55721 59931 55749 59959
rect 55659 59869 55687 59897
rect 55721 59869 55749 59897
rect 55659 59807 55687 59835
rect 55721 59807 55749 59835
rect 55659 59745 55687 59773
rect 55721 59745 55749 59773
rect 71019 59931 71047 59959
rect 71081 59931 71109 59959
rect 71019 59869 71047 59897
rect 71081 59869 71109 59897
rect 71019 59807 71047 59835
rect 71081 59807 71109 59835
rect 71019 59745 71047 59773
rect 71081 59745 71109 59773
rect 86379 59931 86407 59959
rect 86441 59931 86469 59959
rect 86379 59869 86407 59897
rect 86441 59869 86469 59897
rect 86379 59807 86407 59835
rect 86441 59807 86469 59835
rect 86379 59745 86407 59773
rect 86441 59745 86469 59773
rect 101739 59931 101767 59959
rect 101801 59931 101829 59959
rect 101739 59869 101767 59897
rect 101801 59869 101829 59897
rect 101739 59807 101767 59835
rect 101801 59807 101829 59835
rect 101739 59745 101767 59773
rect 101801 59745 101829 59773
rect 117099 59931 117127 59959
rect 117161 59931 117189 59959
rect 117099 59869 117127 59897
rect 117161 59869 117189 59897
rect 117099 59807 117127 59835
rect 117161 59807 117189 59835
rect 117099 59745 117127 59773
rect 117161 59745 117189 59773
rect 132459 59931 132487 59959
rect 132521 59931 132549 59959
rect 132459 59869 132487 59897
rect 132521 59869 132549 59897
rect 132459 59807 132487 59835
rect 132521 59807 132549 59835
rect 132459 59745 132487 59773
rect 132521 59745 132549 59773
rect 147819 59931 147847 59959
rect 147881 59931 147909 59959
rect 147819 59869 147847 59897
rect 147881 59869 147909 59897
rect 147819 59807 147847 59835
rect 147881 59807 147909 59835
rect 147819 59745 147847 59773
rect 147881 59745 147909 59773
rect 163179 59931 163207 59959
rect 163241 59931 163269 59959
rect 163179 59869 163207 59897
rect 163241 59869 163269 59897
rect 163179 59807 163207 59835
rect 163241 59807 163269 59835
rect 163179 59745 163207 59773
rect 163241 59745 163269 59773
rect 178539 59931 178567 59959
rect 178601 59931 178629 59959
rect 178539 59869 178567 59897
rect 178601 59869 178629 59897
rect 178539 59807 178567 59835
rect 178601 59807 178629 59835
rect 178539 59745 178567 59773
rect 178601 59745 178629 59773
rect 193899 59931 193927 59959
rect 193961 59931 193989 59959
rect 193899 59869 193927 59897
rect 193961 59869 193989 59897
rect 193899 59807 193927 59835
rect 193961 59807 193989 59835
rect 193899 59745 193927 59773
rect 193961 59745 193989 59773
rect 209259 59931 209287 59959
rect 209321 59931 209349 59959
rect 209259 59869 209287 59897
rect 209321 59869 209349 59897
rect 209259 59807 209287 59835
rect 209321 59807 209349 59835
rect 209259 59745 209287 59773
rect 209321 59745 209349 59773
rect 224619 59931 224647 59959
rect 224681 59931 224709 59959
rect 224619 59869 224647 59897
rect 224681 59869 224709 59897
rect 224619 59807 224647 59835
rect 224681 59807 224709 59835
rect 224619 59745 224647 59773
rect 224681 59745 224709 59773
rect 239979 59931 240007 59959
rect 240041 59931 240069 59959
rect 239979 59869 240007 59897
rect 240041 59869 240069 59897
rect 239979 59807 240007 59835
rect 240041 59807 240069 59835
rect 239979 59745 240007 59773
rect 240041 59745 240069 59773
rect 32619 56931 32647 56959
rect 32681 56931 32709 56959
rect 32619 56869 32647 56897
rect 32681 56869 32709 56897
rect 32619 56807 32647 56835
rect 32681 56807 32709 56835
rect 32619 56745 32647 56773
rect 32681 56745 32709 56773
rect 47979 56931 48007 56959
rect 48041 56931 48069 56959
rect 47979 56869 48007 56897
rect 48041 56869 48069 56897
rect 47979 56807 48007 56835
rect 48041 56807 48069 56835
rect 47979 56745 48007 56773
rect 48041 56745 48069 56773
rect 63339 56931 63367 56959
rect 63401 56931 63429 56959
rect 63339 56869 63367 56897
rect 63401 56869 63429 56897
rect 63339 56807 63367 56835
rect 63401 56807 63429 56835
rect 63339 56745 63367 56773
rect 63401 56745 63429 56773
rect 78699 56931 78727 56959
rect 78761 56931 78789 56959
rect 78699 56869 78727 56897
rect 78761 56869 78789 56897
rect 78699 56807 78727 56835
rect 78761 56807 78789 56835
rect 78699 56745 78727 56773
rect 78761 56745 78789 56773
rect 94059 56931 94087 56959
rect 94121 56931 94149 56959
rect 94059 56869 94087 56897
rect 94121 56869 94149 56897
rect 94059 56807 94087 56835
rect 94121 56807 94149 56835
rect 94059 56745 94087 56773
rect 94121 56745 94149 56773
rect 109419 56931 109447 56959
rect 109481 56931 109509 56959
rect 109419 56869 109447 56897
rect 109481 56869 109509 56897
rect 109419 56807 109447 56835
rect 109481 56807 109509 56835
rect 109419 56745 109447 56773
rect 109481 56745 109509 56773
rect 124779 56931 124807 56959
rect 124841 56931 124869 56959
rect 124779 56869 124807 56897
rect 124841 56869 124869 56897
rect 124779 56807 124807 56835
rect 124841 56807 124869 56835
rect 124779 56745 124807 56773
rect 124841 56745 124869 56773
rect 140139 56931 140167 56959
rect 140201 56931 140229 56959
rect 140139 56869 140167 56897
rect 140201 56869 140229 56897
rect 140139 56807 140167 56835
rect 140201 56807 140229 56835
rect 140139 56745 140167 56773
rect 140201 56745 140229 56773
rect 155499 56931 155527 56959
rect 155561 56931 155589 56959
rect 155499 56869 155527 56897
rect 155561 56869 155589 56897
rect 155499 56807 155527 56835
rect 155561 56807 155589 56835
rect 155499 56745 155527 56773
rect 155561 56745 155589 56773
rect 170859 56931 170887 56959
rect 170921 56931 170949 56959
rect 170859 56869 170887 56897
rect 170921 56869 170949 56897
rect 170859 56807 170887 56835
rect 170921 56807 170949 56835
rect 170859 56745 170887 56773
rect 170921 56745 170949 56773
rect 186219 56931 186247 56959
rect 186281 56931 186309 56959
rect 186219 56869 186247 56897
rect 186281 56869 186309 56897
rect 186219 56807 186247 56835
rect 186281 56807 186309 56835
rect 186219 56745 186247 56773
rect 186281 56745 186309 56773
rect 201579 56931 201607 56959
rect 201641 56931 201669 56959
rect 201579 56869 201607 56897
rect 201641 56869 201669 56897
rect 201579 56807 201607 56835
rect 201641 56807 201669 56835
rect 201579 56745 201607 56773
rect 201641 56745 201669 56773
rect 216939 56931 216967 56959
rect 217001 56931 217029 56959
rect 216939 56869 216967 56897
rect 217001 56869 217029 56897
rect 216939 56807 216967 56835
rect 217001 56807 217029 56835
rect 216939 56745 216967 56773
rect 217001 56745 217029 56773
rect 232299 56931 232327 56959
rect 232361 56931 232389 56959
rect 232299 56869 232327 56897
rect 232361 56869 232389 56897
rect 232299 56807 232327 56835
rect 232361 56807 232389 56835
rect 232299 56745 232327 56773
rect 232361 56745 232389 56773
rect 247659 56931 247687 56959
rect 247721 56931 247749 56959
rect 247659 56869 247687 56897
rect 247721 56869 247749 56897
rect 247659 56807 247687 56835
rect 247721 56807 247749 56835
rect 247659 56745 247687 56773
rect 247721 56745 247749 56773
rect 254577 56931 254605 56959
rect 254639 56931 254667 56959
rect 254701 56931 254729 56959
rect 254763 56931 254791 56959
rect 254577 56869 254605 56897
rect 254639 56869 254667 56897
rect 254701 56869 254729 56897
rect 254763 56869 254791 56897
rect 254577 56807 254605 56835
rect 254639 56807 254667 56835
rect 254701 56807 254729 56835
rect 254763 56807 254791 56835
rect 254577 56745 254605 56773
rect 254639 56745 254667 56773
rect 254701 56745 254729 56773
rect 254763 56745 254791 56773
rect 31437 50931 31465 50959
rect 31499 50931 31527 50959
rect 31561 50931 31589 50959
rect 31623 50931 31651 50959
rect 31437 50869 31465 50897
rect 31499 50869 31527 50897
rect 31561 50869 31589 50897
rect 31623 50869 31651 50897
rect 31437 50807 31465 50835
rect 31499 50807 31527 50835
rect 31561 50807 31589 50835
rect 31623 50807 31651 50835
rect 31437 50745 31465 50773
rect 31499 50745 31527 50773
rect 31561 50745 31589 50773
rect 31623 50745 31651 50773
rect 40299 50931 40327 50959
rect 40361 50931 40389 50959
rect 40299 50869 40327 50897
rect 40361 50869 40389 50897
rect 40299 50807 40327 50835
rect 40361 50807 40389 50835
rect 40299 50745 40327 50773
rect 40361 50745 40389 50773
rect 55659 50931 55687 50959
rect 55721 50931 55749 50959
rect 55659 50869 55687 50897
rect 55721 50869 55749 50897
rect 55659 50807 55687 50835
rect 55721 50807 55749 50835
rect 55659 50745 55687 50773
rect 55721 50745 55749 50773
rect 71019 50931 71047 50959
rect 71081 50931 71109 50959
rect 71019 50869 71047 50897
rect 71081 50869 71109 50897
rect 71019 50807 71047 50835
rect 71081 50807 71109 50835
rect 71019 50745 71047 50773
rect 71081 50745 71109 50773
rect 86379 50931 86407 50959
rect 86441 50931 86469 50959
rect 86379 50869 86407 50897
rect 86441 50869 86469 50897
rect 86379 50807 86407 50835
rect 86441 50807 86469 50835
rect 86379 50745 86407 50773
rect 86441 50745 86469 50773
rect 101739 50931 101767 50959
rect 101801 50931 101829 50959
rect 101739 50869 101767 50897
rect 101801 50869 101829 50897
rect 101739 50807 101767 50835
rect 101801 50807 101829 50835
rect 101739 50745 101767 50773
rect 101801 50745 101829 50773
rect 117099 50931 117127 50959
rect 117161 50931 117189 50959
rect 117099 50869 117127 50897
rect 117161 50869 117189 50897
rect 117099 50807 117127 50835
rect 117161 50807 117189 50835
rect 117099 50745 117127 50773
rect 117161 50745 117189 50773
rect 132459 50931 132487 50959
rect 132521 50931 132549 50959
rect 132459 50869 132487 50897
rect 132521 50869 132549 50897
rect 132459 50807 132487 50835
rect 132521 50807 132549 50835
rect 132459 50745 132487 50773
rect 132521 50745 132549 50773
rect 147819 50931 147847 50959
rect 147881 50931 147909 50959
rect 147819 50869 147847 50897
rect 147881 50869 147909 50897
rect 147819 50807 147847 50835
rect 147881 50807 147909 50835
rect 147819 50745 147847 50773
rect 147881 50745 147909 50773
rect 163179 50931 163207 50959
rect 163241 50931 163269 50959
rect 163179 50869 163207 50897
rect 163241 50869 163269 50897
rect 163179 50807 163207 50835
rect 163241 50807 163269 50835
rect 163179 50745 163207 50773
rect 163241 50745 163269 50773
rect 178539 50931 178567 50959
rect 178601 50931 178629 50959
rect 178539 50869 178567 50897
rect 178601 50869 178629 50897
rect 178539 50807 178567 50835
rect 178601 50807 178629 50835
rect 178539 50745 178567 50773
rect 178601 50745 178629 50773
rect 193899 50931 193927 50959
rect 193961 50931 193989 50959
rect 193899 50869 193927 50897
rect 193961 50869 193989 50897
rect 193899 50807 193927 50835
rect 193961 50807 193989 50835
rect 193899 50745 193927 50773
rect 193961 50745 193989 50773
rect 209259 50931 209287 50959
rect 209321 50931 209349 50959
rect 209259 50869 209287 50897
rect 209321 50869 209349 50897
rect 209259 50807 209287 50835
rect 209321 50807 209349 50835
rect 209259 50745 209287 50773
rect 209321 50745 209349 50773
rect 224619 50931 224647 50959
rect 224681 50931 224709 50959
rect 224619 50869 224647 50897
rect 224681 50869 224709 50897
rect 224619 50807 224647 50835
rect 224681 50807 224709 50835
rect 224619 50745 224647 50773
rect 224681 50745 224709 50773
rect 239979 50931 240007 50959
rect 240041 50931 240069 50959
rect 239979 50869 240007 50897
rect 240041 50869 240069 50897
rect 239979 50807 240007 50835
rect 240041 50807 240069 50835
rect 239979 50745 240007 50773
rect 240041 50745 240069 50773
rect 32619 47931 32647 47959
rect 32681 47931 32709 47959
rect 32619 47869 32647 47897
rect 32681 47869 32709 47897
rect 32619 47807 32647 47835
rect 32681 47807 32709 47835
rect 32619 47745 32647 47773
rect 32681 47745 32709 47773
rect 47979 47931 48007 47959
rect 48041 47931 48069 47959
rect 47979 47869 48007 47897
rect 48041 47869 48069 47897
rect 47979 47807 48007 47835
rect 48041 47807 48069 47835
rect 47979 47745 48007 47773
rect 48041 47745 48069 47773
rect 63339 47931 63367 47959
rect 63401 47931 63429 47959
rect 63339 47869 63367 47897
rect 63401 47869 63429 47897
rect 63339 47807 63367 47835
rect 63401 47807 63429 47835
rect 63339 47745 63367 47773
rect 63401 47745 63429 47773
rect 78699 47931 78727 47959
rect 78761 47931 78789 47959
rect 78699 47869 78727 47897
rect 78761 47869 78789 47897
rect 78699 47807 78727 47835
rect 78761 47807 78789 47835
rect 78699 47745 78727 47773
rect 78761 47745 78789 47773
rect 94059 47931 94087 47959
rect 94121 47931 94149 47959
rect 94059 47869 94087 47897
rect 94121 47869 94149 47897
rect 94059 47807 94087 47835
rect 94121 47807 94149 47835
rect 94059 47745 94087 47773
rect 94121 47745 94149 47773
rect 109419 47931 109447 47959
rect 109481 47931 109509 47959
rect 109419 47869 109447 47897
rect 109481 47869 109509 47897
rect 109419 47807 109447 47835
rect 109481 47807 109509 47835
rect 109419 47745 109447 47773
rect 109481 47745 109509 47773
rect 124779 47931 124807 47959
rect 124841 47931 124869 47959
rect 124779 47869 124807 47897
rect 124841 47869 124869 47897
rect 124779 47807 124807 47835
rect 124841 47807 124869 47835
rect 124779 47745 124807 47773
rect 124841 47745 124869 47773
rect 140139 47931 140167 47959
rect 140201 47931 140229 47959
rect 140139 47869 140167 47897
rect 140201 47869 140229 47897
rect 140139 47807 140167 47835
rect 140201 47807 140229 47835
rect 140139 47745 140167 47773
rect 140201 47745 140229 47773
rect 155499 47931 155527 47959
rect 155561 47931 155589 47959
rect 155499 47869 155527 47897
rect 155561 47869 155589 47897
rect 155499 47807 155527 47835
rect 155561 47807 155589 47835
rect 155499 47745 155527 47773
rect 155561 47745 155589 47773
rect 170859 47931 170887 47959
rect 170921 47931 170949 47959
rect 170859 47869 170887 47897
rect 170921 47869 170949 47897
rect 170859 47807 170887 47835
rect 170921 47807 170949 47835
rect 170859 47745 170887 47773
rect 170921 47745 170949 47773
rect 186219 47931 186247 47959
rect 186281 47931 186309 47959
rect 186219 47869 186247 47897
rect 186281 47869 186309 47897
rect 186219 47807 186247 47835
rect 186281 47807 186309 47835
rect 186219 47745 186247 47773
rect 186281 47745 186309 47773
rect 201579 47931 201607 47959
rect 201641 47931 201669 47959
rect 201579 47869 201607 47897
rect 201641 47869 201669 47897
rect 201579 47807 201607 47835
rect 201641 47807 201669 47835
rect 201579 47745 201607 47773
rect 201641 47745 201669 47773
rect 216939 47931 216967 47959
rect 217001 47931 217029 47959
rect 216939 47869 216967 47897
rect 217001 47869 217029 47897
rect 216939 47807 216967 47835
rect 217001 47807 217029 47835
rect 216939 47745 216967 47773
rect 217001 47745 217029 47773
rect 232299 47931 232327 47959
rect 232361 47931 232389 47959
rect 232299 47869 232327 47897
rect 232361 47869 232389 47897
rect 232299 47807 232327 47835
rect 232361 47807 232389 47835
rect 232299 47745 232327 47773
rect 232361 47745 232389 47773
rect 247659 47931 247687 47959
rect 247721 47931 247749 47959
rect 247659 47869 247687 47897
rect 247721 47869 247749 47897
rect 247659 47807 247687 47835
rect 247721 47807 247749 47835
rect 247659 47745 247687 47773
rect 247721 47745 247749 47773
rect 254577 47931 254605 47959
rect 254639 47931 254667 47959
rect 254701 47931 254729 47959
rect 254763 47931 254791 47959
rect 254577 47869 254605 47897
rect 254639 47869 254667 47897
rect 254701 47869 254729 47897
rect 254763 47869 254791 47897
rect 254577 47807 254605 47835
rect 254639 47807 254667 47835
rect 254701 47807 254729 47835
rect 254763 47807 254791 47835
rect 254577 47745 254605 47773
rect 254639 47745 254667 47773
rect 254701 47745 254729 47773
rect 254763 47745 254791 47773
rect 31437 41931 31465 41959
rect 31499 41931 31527 41959
rect 31561 41931 31589 41959
rect 31623 41931 31651 41959
rect 31437 41869 31465 41897
rect 31499 41869 31527 41897
rect 31561 41869 31589 41897
rect 31623 41869 31651 41897
rect 31437 41807 31465 41835
rect 31499 41807 31527 41835
rect 31561 41807 31589 41835
rect 31623 41807 31651 41835
rect 31437 41745 31465 41773
rect 31499 41745 31527 41773
rect 31561 41745 31589 41773
rect 31623 41745 31651 41773
rect 40299 41931 40327 41959
rect 40361 41931 40389 41959
rect 40299 41869 40327 41897
rect 40361 41869 40389 41897
rect 40299 41807 40327 41835
rect 40361 41807 40389 41835
rect 40299 41745 40327 41773
rect 40361 41745 40389 41773
rect 55659 41931 55687 41959
rect 55721 41931 55749 41959
rect 55659 41869 55687 41897
rect 55721 41869 55749 41897
rect 55659 41807 55687 41835
rect 55721 41807 55749 41835
rect 55659 41745 55687 41773
rect 55721 41745 55749 41773
rect 71019 41931 71047 41959
rect 71081 41931 71109 41959
rect 71019 41869 71047 41897
rect 71081 41869 71109 41897
rect 71019 41807 71047 41835
rect 71081 41807 71109 41835
rect 71019 41745 71047 41773
rect 71081 41745 71109 41773
rect 86379 41931 86407 41959
rect 86441 41931 86469 41959
rect 86379 41869 86407 41897
rect 86441 41869 86469 41897
rect 86379 41807 86407 41835
rect 86441 41807 86469 41835
rect 86379 41745 86407 41773
rect 86441 41745 86469 41773
rect 101739 41931 101767 41959
rect 101801 41931 101829 41959
rect 101739 41869 101767 41897
rect 101801 41869 101829 41897
rect 101739 41807 101767 41835
rect 101801 41807 101829 41835
rect 101739 41745 101767 41773
rect 101801 41745 101829 41773
rect 117099 41931 117127 41959
rect 117161 41931 117189 41959
rect 117099 41869 117127 41897
rect 117161 41869 117189 41897
rect 117099 41807 117127 41835
rect 117161 41807 117189 41835
rect 117099 41745 117127 41773
rect 117161 41745 117189 41773
rect 132459 41931 132487 41959
rect 132521 41931 132549 41959
rect 132459 41869 132487 41897
rect 132521 41869 132549 41897
rect 132459 41807 132487 41835
rect 132521 41807 132549 41835
rect 132459 41745 132487 41773
rect 132521 41745 132549 41773
rect 147819 41931 147847 41959
rect 147881 41931 147909 41959
rect 147819 41869 147847 41897
rect 147881 41869 147909 41897
rect 147819 41807 147847 41835
rect 147881 41807 147909 41835
rect 147819 41745 147847 41773
rect 147881 41745 147909 41773
rect 163179 41931 163207 41959
rect 163241 41931 163269 41959
rect 163179 41869 163207 41897
rect 163241 41869 163269 41897
rect 163179 41807 163207 41835
rect 163241 41807 163269 41835
rect 163179 41745 163207 41773
rect 163241 41745 163269 41773
rect 178539 41931 178567 41959
rect 178601 41931 178629 41959
rect 178539 41869 178567 41897
rect 178601 41869 178629 41897
rect 178539 41807 178567 41835
rect 178601 41807 178629 41835
rect 178539 41745 178567 41773
rect 178601 41745 178629 41773
rect 193899 41931 193927 41959
rect 193961 41931 193989 41959
rect 193899 41869 193927 41897
rect 193961 41869 193989 41897
rect 193899 41807 193927 41835
rect 193961 41807 193989 41835
rect 193899 41745 193927 41773
rect 193961 41745 193989 41773
rect 209259 41931 209287 41959
rect 209321 41931 209349 41959
rect 209259 41869 209287 41897
rect 209321 41869 209349 41897
rect 209259 41807 209287 41835
rect 209321 41807 209349 41835
rect 209259 41745 209287 41773
rect 209321 41745 209349 41773
rect 224619 41931 224647 41959
rect 224681 41931 224709 41959
rect 224619 41869 224647 41897
rect 224681 41869 224709 41897
rect 224619 41807 224647 41835
rect 224681 41807 224709 41835
rect 224619 41745 224647 41773
rect 224681 41745 224709 41773
rect 239979 41931 240007 41959
rect 240041 41931 240069 41959
rect 239979 41869 240007 41897
rect 240041 41869 240069 41897
rect 239979 41807 240007 41835
rect 240041 41807 240069 41835
rect 239979 41745 240007 41773
rect 240041 41745 240069 41773
rect 32619 38931 32647 38959
rect 32681 38931 32709 38959
rect 32619 38869 32647 38897
rect 32681 38869 32709 38897
rect 32619 38807 32647 38835
rect 32681 38807 32709 38835
rect 32619 38745 32647 38773
rect 32681 38745 32709 38773
rect 47979 38931 48007 38959
rect 48041 38931 48069 38959
rect 47979 38869 48007 38897
rect 48041 38869 48069 38897
rect 47979 38807 48007 38835
rect 48041 38807 48069 38835
rect 47979 38745 48007 38773
rect 48041 38745 48069 38773
rect 63339 38931 63367 38959
rect 63401 38931 63429 38959
rect 63339 38869 63367 38897
rect 63401 38869 63429 38897
rect 63339 38807 63367 38835
rect 63401 38807 63429 38835
rect 63339 38745 63367 38773
rect 63401 38745 63429 38773
rect 78699 38931 78727 38959
rect 78761 38931 78789 38959
rect 78699 38869 78727 38897
rect 78761 38869 78789 38897
rect 78699 38807 78727 38835
rect 78761 38807 78789 38835
rect 78699 38745 78727 38773
rect 78761 38745 78789 38773
rect 94059 38931 94087 38959
rect 94121 38931 94149 38959
rect 94059 38869 94087 38897
rect 94121 38869 94149 38897
rect 94059 38807 94087 38835
rect 94121 38807 94149 38835
rect 94059 38745 94087 38773
rect 94121 38745 94149 38773
rect 109419 38931 109447 38959
rect 109481 38931 109509 38959
rect 109419 38869 109447 38897
rect 109481 38869 109509 38897
rect 109419 38807 109447 38835
rect 109481 38807 109509 38835
rect 109419 38745 109447 38773
rect 109481 38745 109509 38773
rect 124779 38931 124807 38959
rect 124841 38931 124869 38959
rect 124779 38869 124807 38897
rect 124841 38869 124869 38897
rect 124779 38807 124807 38835
rect 124841 38807 124869 38835
rect 124779 38745 124807 38773
rect 124841 38745 124869 38773
rect 140139 38931 140167 38959
rect 140201 38931 140229 38959
rect 140139 38869 140167 38897
rect 140201 38869 140229 38897
rect 140139 38807 140167 38835
rect 140201 38807 140229 38835
rect 140139 38745 140167 38773
rect 140201 38745 140229 38773
rect 155499 38931 155527 38959
rect 155561 38931 155589 38959
rect 155499 38869 155527 38897
rect 155561 38869 155589 38897
rect 155499 38807 155527 38835
rect 155561 38807 155589 38835
rect 155499 38745 155527 38773
rect 155561 38745 155589 38773
rect 170859 38931 170887 38959
rect 170921 38931 170949 38959
rect 170859 38869 170887 38897
rect 170921 38869 170949 38897
rect 170859 38807 170887 38835
rect 170921 38807 170949 38835
rect 170859 38745 170887 38773
rect 170921 38745 170949 38773
rect 186219 38931 186247 38959
rect 186281 38931 186309 38959
rect 186219 38869 186247 38897
rect 186281 38869 186309 38897
rect 186219 38807 186247 38835
rect 186281 38807 186309 38835
rect 186219 38745 186247 38773
rect 186281 38745 186309 38773
rect 201579 38931 201607 38959
rect 201641 38931 201669 38959
rect 201579 38869 201607 38897
rect 201641 38869 201669 38897
rect 201579 38807 201607 38835
rect 201641 38807 201669 38835
rect 201579 38745 201607 38773
rect 201641 38745 201669 38773
rect 216939 38931 216967 38959
rect 217001 38931 217029 38959
rect 216939 38869 216967 38897
rect 217001 38869 217029 38897
rect 216939 38807 216967 38835
rect 217001 38807 217029 38835
rect 216939 38745 216967 38773
rect 217001 38745 217029 38773
rect 232299 38931 232327 38959
rect 232361 38931 232389 38959
rect 232299 38869 232327 38897
rect 232361 38869 232389 38897
rect 232299 38807 232327 38835
rect 232361 38807 232389 38835
rect 232299 38745 232327 38773
rect 232361 38745 232389 38773
rect 247659 38931 247687 38959
rect 247721 38931 247749 38959
rect 247659 38869 247687 38897
rect 247721 38869 247749 38897
rect 247659 38807 247687 38835
rect 247721 38807 247749 38835
rect 247659 38745 247687 38773
rect 247721 38745 247749 38773
rect 254577 38931 254605 38959
rect 254639 38931 254667 38959
rect 254701 38931 254729 38959
rect 254763 38931 254791 38959
rect 254577 38869 254605 38897
rect 254639 38869 254667 38897
rect 254701 38869 254729 38897
rect 254763 38869 254791 38897
rect 254577 38807 254605 38835
rect 254639 38807 254667 38835
rect 254701 38807 254729 38835
rect 254763 38807 254791 38835
rect 254577 38745 254605 38773
rect 254639 38745 254667 38773
rect 254701 38745 254729 38773
rect 254763 38745 254791 38773
rect 31437 32931 31465 32959
rect 31499 32931 31527 32959
rect 31561 32931 31589 32959
rect 31623 32931 31651 32959
rect 31437 32869 31465 32897
rect 31499 32869 31527 32897
rect 31561 32869 31589 32897
rect 31623 32869 31651 32897
rect 31437 32807 31465 32835
rect 31499 32807 31527 32835
rect 31561 32807 31589 32835
rect 31623 32807 31651 32835
rect 31437 32745 31465 32773
rect 31499 32745 31527 32773
rect 31561 32745 31589 32773
rect 31623 32745 31651 32773
rect 40299 32931 40327 32959
rect 40361 32931 40389 32959
rect 40299 32869 40327 32897
rect 40361 32869 40389 32897
rect 40299 32807 40327 32835
rect 40361 32807 40389 32835
rect 40299 32745 40327 32773
rect 40361 32745 40389 32773
rect 55659 32931 55687 32959
rect 55721 32931 55749 32959
rect 55659 32869 55687 32897
rect 55721 32869 55749 32897
rect 55659 32807 55687 32835
rect 55721 32807 55749 32835
rect 55659 32745 55687 32773
rect 55721 32745 55749 32773
rect 71019 32931 71047 32959
rect 71081 32931 71109 32959
rect 71019 32869 71047 32897
rect 71081 32869 71109 32897
rect 71019 32807 71047 32835
rect 71081 32807 71109 32835
rect 71019 32745 71047 32773
rect 71081 32745 71109 32773
rect 86379 32931 86407 32959
rect 86441 32931 86469 32959
rect 86379 32869 86407 32897
rect 86441 32869 86469 32897
rect 86379 32807 86407 32835
rect 86441 32807 86469 32835
rect 86379 32745 86407 32773
rect 86441 32745 86469 32773
rect 101739 32931 101767 32959
rect 101801 32931 101829 32959
rect 101739 32869 101767 32897
rect 101801 32869 101829 32897
rect 101739 32807 101767 32835
rect 101801 32807 101829 32835
rect 101739 32745 101767 32773
rect 101801 32745 101829 32773
rect 117099 32931 117127 32959
rect 117161 32931 117189 32959
rect 117099 32869 117127 32897
rect 117161 32869 117189 32897
rect 117099 32807 117127 32835
rect 117161 32807 117189 32835
rect 117099 32745 117127 32773
rect 117161 32745 117189 32773
rect 132459 32931 132487 32959
rect 132521 32931 132549 32959
rect 132459 32869 132487 32897
rect 132521 32869 132549 32897
rect 132459 32807 132487 32835
rect 132521 32807 132549 32835
rect 132459 32745 132487 32773
rect 132521 32745 132549 32773
rect 147819 32931 147847 32959
rect 147881 32931 147909 32959
rect 147819 32869 147847 32897
rect 147881 32869 147909 32897
rect 147819 32807 147847 32835
rect 147881 32807 147909 32835
rect 147819 32745 147847 32773
rect 147881 32745 147909 32773
rect 163179 32931 163207 32959
rect 163241 32931 163269 32959
rect 163179 32869 163207 32897
rect 163241 32869 163269 32897
rect 163179 32807 163207 32835
rect 163241 32807 163269 32835
rect 163179 32745 163207 32773
rect 163241 32745 163269 32773
rect 178539 32931 178567 32959
rect 178601 32931 178629 32959
rect 178539 32869 178567 32897
rect 178601 32869 178629 32897
rect 178539 32807 178567 32835
rect 178601 32807 178629 32835
rect 178539 32745 178567 32773
rect 178601 32745 178629 32773
rect 193899 32931 193927 32959
rect 193961 32931 193989 32959
rect 193899 32869 193927 32897
rect 193961 32869 193989 32897
rect 193899 32807 193927 32835
rect 193961 32807 193989 32835
rect 193899 32745 193927 32773
rect 193961 32745 193989 32773
rect 209259 32931 209287 32959
rect 209321 32931 209349 32959
rect 209259 32869 209287 32897
rect 209321 32869 209349 32897
rect 209259 32807 209287 32835
rect 209321 32807 209349 32835
rect 209259 32745 209287 32773
rect 209321 32745 209349 32773
rect 224619 32931 224647 32959
rect 224681 32931 224709 32959
rect 224619 32869 224647 32897
rect 224681 32869 224709 32897
rect 224619 32807 224647 32835
rect 224681 32807 224709 32835
rect 224619 32745 224647 32773
rect 224681 32745 224709 32773
rect 239979 32931 240007 32959
rect 240041 32931 240069 32959
rect 239979 32869 240007 32897
rect 240041 32869 240069 32897
rect 239979 32807 240007 32835
rect 240041 32807 240069 32835
rect 239979 32745 240007 32773
rect 240041 32745 240069 32773
rect 32619 29931 32647 29959
rect 32681 29931 32709 29959
rect 32619 29869 32647 29897
rect 32681 29869 32709 29897
rect 32619 29807 32647 29835
rect 32681 29807 32709 29835
rect 32619 29745 32647 29773
rect 32681 29745 32709 29773
rect 47979 29931 48007 29959
rect 48041 29931 48069 29959
rect 47979 29869 48007 29897
rect 48041 29869 48069 29897
rect 47979 29807 48007 29835
rect 48041 29807 48069 29835
rect 47979 29745 48007 29773
rect 48041 29745 48069 29773
rect 63339 29931 63367 29959
rect 63401 29931 63429 29959
rect 63339 29869 63367 29897
rect 63401 29869 63429 29897
rect 63339 29807 63367 29835
rect 63401 29807 63429 29835
rect 63339 29745 63367 29773
rect 63401 29745 63429 29773
rect 78699 29931 78727 29959
rect 78761 29931 78789 29959
rect 78699 29869 78727 29897
rect 78761 29869 78789 29897
rect 78699 29807 78727 29835
rect 78761 29807 78789 29835
rect 78699 29745 78727 29773
rect 78761 29745 78789 29773
rect 94059 29931 94087 29959
rect 94121 29931 94149 29959
rect 94059 29869 94087 29897
rect 94121 29869 94149 29897
rect 94059 29807 94087 29835
rect 94121 29807 94149 29835
rect 94059 29745 94087 29773
rect 94121 29745 94149 29773
rect 109419 29931 109447 29959
rect 109481 29931 109509 29959
rect 109419 29869 109447 29897
rect 109481 29869 109509 29897
rect 109419 29807 109447 29835
rect 109481 29807 109509 29835
rect 109419 29745 109447 29773
rect 109481 29745 109509 29773
rect 124779 29931 124807 29959
rect 124841 29931 124869 29959
rect 124779 29869 124807 29897
rect 124841 29869 124869 29897
rect 124779 29807 124807 29835
rect 124841 29807 124869 29835
rect 124779 29745 124807 29773
rect 124841 29745 124869 29773
rect 140139 29931 140167 29959
rect 140201 29931 140229 29959
rect 140139 29869 140167 29897
rect 140201 29869 140229 29897
rect 140139 29807 140167 29835
rect 140201 29807 140229 29835
rect 140139 29745 140167 29773
rect 140201 29745 140229 29773
rect 155499 29931 155527 29959
rect 155561 29931 155589 29959
rect 155499 29869 155527 29897
rect 155561 29869 155589 29897
rect 155499 29807 155527 29835
rect 155561 29807 155589 29835
rect 155499 29745 155527 29773
rect 155561 29745 155589 29773
rect 170859 29931 170887 29959
rect 170921 29931 170949 29959
rect 170859 29869 170887 29897
rect 170921 29869 170949 29897
rect 170859 29807 170887 29835
rect 170921 29807 170949 29835
rect 170859 29745 170887 29773
rect 170921 29745 170949 29773
rect 186219 29931 186247 29959
rect 186281 29931 186309 29959
rect 186219 29869 186247 29897
rect 186281 29869 186309 29897
rect 186219 29807 186247 29835
rect 186281 29807 186309 29835
rect 186219 29745 186247 29773
rect 186281 29745 186309 29773
rect 201579 29931 201607 29959
rect 201641 29931 201669 29959
rect 201579 29869 201607 29897
rect 201641 29869 201669 29897
rect 201579 29807 201607 29835
rect 201641 29807 201669 29835
rect 201579 29745 201607 29773
rect 201641 29745 201669 29773
rect 216939 29931 216967 29959
rect 217001 29931 217029 29959
rect 216939 29869 216967 29897
rect 217001 29869 217029 29897
rect 216939 29807 216967 29835
rect 217001 29807 217029 29835
rect 216939 29745 216967 29773
rect 217001 29745 217029 29773
rect 232299 29931 232327 29959
rect 232361 29931 232389 29959
rect 232299 29869 232327 29897
rect 232361 29869 232389 29897
rect 232299 29807 232327 29835
rect 232361 29807 232389 29835
rect 232299 29745 232327 29773
rect 232361 29745 232389 29773
rect 247659 29931 247687 29959
rect 247721 29931 247749 29959
rect 247659 29869 247687 29897
rect 247721 29869 247749 29897
rect 247659 29807 247687 29835
rect 247721 29807 247749 29835
rect 247659 29745 247687 29773
rect 247721 29745 247749 29773
rect 254577 29931 254605 29959
rect 254639 29931 254667 29959
rect 254701 29931 254729 29959
rect 254763 29931 254791 29959
rect 254577 29869 254605 29897
rect 254639 29869 254667 29897
rect 254701 29869 254729 29897
rect 254763 29869 254791 29897
rect 254577 29807 254605 29835
rect 254639 29807 254667 29835
rect 254701 29807 254729 29835
rect 254763 29807 254791 29835
rect 254577 29745 254605 29773
rect 254639 29745 254667 29773
rect 254701 29745 254729 29773
rect 254763 29745 254791 29773
rect 31437 23931 31465 23959
rect 31499 23931 31527 23959
rect 31561 23931 31589 23959
rect 31623 23931 31651 23959
rect 31437 23869 31465 23897
rect 31499 23869 31527 23897
rect 31561 23869 31589 23897
rect 31623 23869 31651 23897
rect 31437 23807 31465 23835
rect 31499 23807 31527 23835
rect 31561 23807 31589 23835
rect 31623 23807 31651 23835
rect 31437 23745 31465 23773
rect 31499 23745 31527 23773
rect 31561 23745 31589 23773
rect 31623 23745 31651 23773
rect 40299 23931 40327 23959
rect 40361 23931 40389 23959
rect 40299 23869 40327 23897
rect 40361 23869 40389 23897
rect 40299 23807 40327 23835
rect 40361 23807 40389 23835
rect 40299 23745 40327 23773
rect 40361 23745 40389 23773
rect 55659 23931 55687 23959
rect 55721 23931 55749 23959
rect 55659 23869 55687 23897
rect 55721 23869 55749 23897
rect 55659 23807 55687 23835
rect 55721 23807 55749 23835
rect 55659 23745 55687 23773
rect 55721 23745 55749 23773
rect 71019 23931 71047 23959
rect 71081 23931 71109 23959
rect 71019 23869 71047 23897
rect 71081 23869 71109 23897
rect 71019 23807 71047 23835
rect 71081 23807 71109 23835
rect 71019 23745 71047 23773
rect 71081 23745 71109 23773
rect 86379 23931 86407 23959
rect 86441 23931 86469 23959
rect 86379 23869 86407 23897
rect 86441 23869 86469 23897
rect 86379 23807 86407 23835
rect 86441 23807 86469 23835
rect 86379 23745 86407 23773
rect 86441 23745 86469 23773
rect 101739 23931 101767 23959
rect 101801 23931 101829 23959
rect 101739 23869 101767 23897
rect 101801 23869 101829 23897
rect 101739 23807 101767 23835
rect 101801 23807 101829 23835
rect 101739 23745 101767 23773
rect 101801 23745 101829 23773
rect 117099 23931 117127 23959
rect 117161 23931 117189 23959
rect 117099 23869 117127 23897
rect 117161 23869 117189 23897
rect 117099 23807 117127 23835
rect 117161 23807 117189 23835
rect 117099 23745 117127 23773
rect 117161 23745 117189 23773
rect 132459 23931 132487 23959
rect 132521 23931 132549 23959
rect 132459 23869 132487 23897
rect 132521 23869 132549 23897
rect 132459 23807 132487 23835
rect 132521 23807 132549 23835
rect 132459 23745 132487 23773
rect 132521 23745 132549 23773
rect 147819 23931 147847 23959
rect 147881 23931 147909 23959
rect 147819 23869 147847 23897
rect 147881 23869 147909 23897
rect 147819 23807 147847 23835
rect 147881 23807 147909 23835
rect 147819 23745 147847 23773
rect 147881 23745 147909 23773
rect 163179 23931 163207 23959
rect 163241 23931 163269 23959
rect 163179 23869 163207 23897
rect 163241 23869 163269 23897
rect 163179 23807 163207 23835
rect 163241 23807 163269 23835
rect 163179 23745 163207 23773
rect 163241 23745 163269 23773
rect 178539 23931 178567 23959
rect 178601 23931 178629 23959
rect 178539 23869 178567 23897
rect 178601 23869 178629 23897
rect 178539 23807 178567 23835
rect 178601 23807 178629 23835
rect 178539 23745 178567 23773
rect 178601 23745 178629 23773
rect 193899 23931 193927 23959
rect 193961 23931 193989 23959
rect 193899 23869 193927 23897
rect 193961 23869 193989 23897
rect 193899 23807 193927 23835
rect 193961 23807 193989 23835
rect 193899 23745 193927 23773
rect 193961 23745 193989 23773
rect 209259 23931 209287 23959
rect 209321 23931 209349 23959
rect 209259 23869 209287 23897
rect 209321 23869 209349 23897
rect 209259 23807 209287 23835
rect 209321 23807 209349 23835
rect 209259 23745 209287 23773
rect 209321 23745 209349 23773
rect 224619 23931 224647 23959
rect 224681 23931 224709 23959
rect 224619 23869 224647 23897
rect 224681 23869 224709 23897
rect 224619 23807 224647 23835
rect 224681 23807 224709 23835
rect 224619 23745 224647 23773
rect 224681 23745 224709 23773
rect 239979 23931 240007 23959
rect 240041 23931 240069 23959
rect 239979 23869 240007 23897
rect 240041 23869 240069 23897
rect 239979 23807 240007 23835
rect 240041 23807 240069 23835
rect 239979 23745 240007 23773
rect 240041 23745 240069 23773
rect 32619 20931 32647 20959
rect 32681 20931 32709 20959
rect 32619 20869 32647 20897
rect 32681 20869 32709 20897
rect 32619 20807 32647 20835
rect 32681 20807 32709 20835
rect 32619 20745 32647 20773
rect 32681 20745 32709 20773
rect 47979 20931 48007 20959
rect 48041 20931 48069 20959
rect 47979 20869 48007 20897
rect 48041 20869 48069 20897
rect 47979 20807 48007 20835
rect 48041 20807 48069 20835
rect 47979 20745 48007 20773
rect 48041 20745 48069 20773
rect 63339 20931 63367 20959
rect 63401 20931 63429 20959
rect 63339 20869 63367 20897
rect 63401 20869 63429 20897
rect 63339 20807 63367 20835
rect 63401 20807 63429 20835
rect 63339 20745 63367 20773
rect 63401 20745 63429 20773
rect 78699 20931 78727 20959
rect 78761 20931 78789 20959
rect 78699 20869 78727 20897
rect 78761 20869 78789 20897
rect 78699 20807 78727 20835
rect 78761 20807 78789 20835
rect 78699 20745 78727 20773
rect 78761 20745 78789 20773
rect 94059 20931 94087 20959
rect 94121 20931 94149 20959
rect 94059 20869 94087 20897
rect 94121 20869 94149 20897
rect 94059 20807 94087 20835
rect 94121 20807 94149 20835
rect 94059 20745 94087 20773
rect 94121 20745 94149 20773
rect 109419 20931 109447 20959
rect 109481 20931 109509 20959
rect 109419 20869 109447 20897
rect 109481 20869 109509 20897
rect 109419 20807 109447 20835
rect 109481 20807 109509 20835
rect 109419 20745 109447 20773
rect 109481 20745 109509 20773
rect 124779 20931 124807 20959
rect 124841 20931 124869 20959
rect 124779 20869 124807 20897
rect 124841 20869 124869 20897
rect 124779 20807 124807 20835
rect 124841 20807 124869 20835
rect 124779 20745 124807 20773
rect 124841 20745 124869 20773
rect 140139 20931 140167 20959
rect 140201 20931 140229 20959
rect 140139 20869 140167 20897
rect 140201 20869 140229 20897
rect 140139 20807 140167 20835
rect 140201 20807 140229 20835
rect 140139 20745 140167 20773
rect 140201 20745 140229 20773
rect 155499 20931 155527 20959
rect 155561 20931 155589 20959
rect 155499 20869 155527 20897
rect 155561 20869 155589 20897
rect 155499 20807 155527 20835
rect 155561 20807 155589 20835
rect 155499 20745 155527 20773
rect 155561 20745 155589 20773
rect 170859 20931 170887 20959
rect 170921 20931 170949 20959
rect 170859 20869 170887 20897
rect 170921 20869 170949 20897
rect 170859 20807 170887 20835
rect 170921 20807 170949 20835
rect 170859 20745 170887 20773
rect 170921 20745 170949 20773
rect 186219 20931 186247 20959
rect 186281 20931 186309 20959
rect 186219 20869 186247 20897
rect 186281 20869 186309 20897
rect 186219 20807 186247 20835
rect 186281 20807 186309 20835
rect 186219 20745 186247 20773
rect 186281 20745 186309 20773
rect 201579 20931 201607 20959
rect 201641 20931 201669 20959
rect 201579 20869 201607 20897
rect 201641 20869 201669 20897
rect 201579 20807 201607 20835
rect 201641 20807 201669 20835
rect 201579 20745 201607 20773
rect 201641 20745 201669 20773
rect 216939 20931 216967 20959
rect 217001 20931 217029 20959
rect 216939 20869 216967 20897
rect 217001 20869 217029 20897
rect 216939 20807 216967 20835
rect 217001 20807 217029 20835
rect 216939 20745 216967 20773
rect 217001 20745 217029 20773
rect 232299 20931 232327 20959
rect 232361 20931 232389 20959
rect 232299 20869 232327 20897
rect 232361 20869 232389 20897
rect 232299 20807 232327 20835
rect 232361 20807 232389 20835
rect 232299 20745 232327 20773
rect 232361 20745 232389 20773
rect 247659 20931 247687 20959
rect 247721 20931 247749 20959
rect 247659 20869 247687 20897
rect 247721 20869 247749 20897
rect 247659 20807 247687 20835
rect 247721 20807 247749 20835
rect 247659 20745 247687 20773
rect 247721 20745 247749 20773
rect 254577 20931 254605 20959
rect 254639 20931 254667 20959
rect 254701 20931 254729 20959
rect 254763 20931 254791 20959
rect 254577 20869 254605 20897
rect 254639 20869 254667 20897
rect 254701 20869 254729 20897
rect 254763 20869 254791 20897
rect 254577 20807 254605 20835
rect 254639 20807 254667 20835
rect 254701 20807 254729 20835
rect 254763 20807 254791 20835
rect 254577 20745 254605 20773
rect 254639 20745 254667 20773
rect 254701 20745 254729 20773
rect 254763 20745 254791 20773
rect 31437 14931 31465 14959
rect 31499 14931 31527 14959
rect 31561 14931 31589 14959
rect 31623 14931 31651 14959
rect 31437 14869 31465 14897
rect 31499 14869 31527 14897
rect 31561 14869 31589 14897
rect 31623 14869 31651 14897
rect 31437 14807 31465 14835
rect 31499 14807 31527 14835
rect 31561 14807 31589 14835
rect 31623 14807 31651 14835
rect 31437 14745 31465 14773
rect 31499 14745 31527 14773
rect 31561 14745 31589 14773
rect 31623 14745 31651 14773
rect 247437 14931 247465 14959
rect 247499 14931 247527 14959
rect 247561 14931 247589 14959
rect 247623 14931 247651 14959
rect 247437 14869 247465 14897
rect 247499 14869 247527 14897
rect 247561 14869 247589 14897
rect 247623 14869 247651 14897
rect 247437 14807 247465 14835
rect 247499 14807 247527 14835
rect 247561 14807 247589 14835
rect 247623 14807 247651 14835
rect 247437 14745 247465 14773
rect 247499 14745 247527 14773
rect 247561 14745 247589 14773
rect 247623 14745 247651 14773
rect 31437 5931 31465 5959
rect 31499 5931 31527 5959
rect 31561 5931 31589 5959
rect 31623 5931 31651 5959
rect 31437 5869 31465 5897
rect 31499 5869 31527 5897
rect 31561 5869 31589 5897
rect 31623 5869 31651 5897
rect 31437 5807 31465 5835
rect 31499 5807 31527 5835
rect 31561 5807 31589 5835
rect 31623 5807 31651 5835
rect 31437 5745 31465 5773
rect 31499 5745 31527 5773
rect 31561 5745 31589 5773
rect 31623 5745 31651 5773
rect 31437 396 31465 424
rect 31499 396 31527 424
rect 31561 396 31589 424
rect 31623 396 31651 424
rect 31437 334 31465 362
rect 31499 334 31527 362
rect 31561 334 31589 362
rect 31623 334 31651 362
rect 31437 272 31465 300
rect 31499 272 31527 300
rect 31561 272 31589 300
rect 31623 272 31651 300
rect 31437 210 31465 238
rect 31499 210 31527 238
rect 31561 210 31589 238
rect 31623 210 31651 238
rect 38577 11931 38605 11959
rect 38639 11931 38667 11959
rect 38701 11931 38729 11959
rect 38763 11931 38791 11959
rect 38577 11869 38605 11897
rect 38639 11869 38667 11897
rect 38701 11869 38729 11897
rect 38763 11869 38791 11897
rect 38577 11807 38605 11835
rect 38639 11807 38667 11835
rect 38701 11807 38729 11835
rect 38763 11807 38791 11835
rect 38577 11745 38605 11773
rect 38639 11745 38667 11773
rect 38701 11745 38729 11773
rect 38763 11745 38791 11773
rect 38577 2931 38605 2959
rect 38639 2931 38667 2959
rect 38701 2931 38729 2959
rect 38763 2931 38791 2959
rect 38577 2869 38605 2897
rect 38639 2869 38667 2897
rect 38701 2869 38729 2897
rect 38763 2869 38791 2897
rect 38577 2807 38605 2835
rect 38639 2807 38667 2835
rect 38701 2807 38729 2835
rect 38763 2807 38791 2835
rect 38577 2745 38605 2773
rect 38639 2745 38667 2773
rect 38701 2745 38729 2773
rect 38763 2745 38791 2773
rect 38577 876 38605 904
rect 38639 876 38667 904
rect 38701 876 38729 904
rect 38763 876 38791 904
rect 38577 814 38605 842
rect 38639 814 38667 842
rect 38701 814 38729 842
rect 38763 814 38791 842
rect 38577 752 38605 780
rect 38639 752 38667 780
rect 38701 752 38729 780
rect 38763 752 38791 780
rect 38577 690 38605 718
rect 38639 690 38667 718
rect 38701 690 38729 718
rect 38763 690 38791 718
rect 40437 5931 40465 5959
rect 40499 5931 40527 5959
rect 40561 5931 40589 5959
rect 40623 5931 40651 5959
rect 40437 5869 40465 5897
rect 40499 5869 40527 5897
rect 40561 5869 40589 5897
rect 40623 5869 40651 5897
rect 40437 5807 40465 5835
rect 40499 5807 40527 5835
rect 40561 5807 40589 5835
rect 40623 5807 40651 5835
rect 40437 5745 40465 5773
rect 40499 5745 40527 5773
rect 40561 5745 40589 5773
rect 40623 5745 40651 5773
rect 40437 396 40465 424
rect 40499 396 40527 424
rect 40561 396 40589 424
rect 40623 396 40651 424
rect 40437 334 40465 362
rect 40499 334 40527 362
rect 40561 334 40589 362
rect 40623 334 40651 362
rect 40437 272 40465 300
rect 40499 272 40527 300
rect 40561 272 40589 300
rect 40623 272 40651 300
rect 40437 210 40465 238
rect 40499 210 40527 238
rect 40561 210 40589 238
rect 40623 210 40651 238
rect 47577 11931 47605 11959
rect 47639 11931 47667 11959
rect 47701 11931 47729 11959
rect 47763 11931 47791 11959
rect 47577 11869 47605 11897
rect 47639 11869 47667 11897
rect 47701 11869 47729 11897
rect 47763 11869 47791 11897
rect 47577 11807 47605 11835
rect 47639 11807 47667 11835
rect 47701 11807 47729 11835
rect 47763 11807 47791 11835
rect 47577 11745 47605 11773
rect 47639 11745 47667 11773
rect 47701 11745 47729 11773
rect 47763 11745 47791 11773
rect 47577 2931 47605 2959
rect 47639 2931 47667 2959
rect 47701 2931 47729 2959
rect 47763 2931 47791 2959
rect 47577 2869 47605 2897
rect 47639 2869 47667 2897
rect 47701 2869 47729 2897
rect 47763 2869 47791 2897
rect 47577 2807 47605 2835
rect 47639 2807 47667 2835
rect 47701 2807 47729 2835
rect 47763 2807 47791 2835
rect 47577 2745 47605 2773
rect 47639 2745 47667 2773
rect 47701 2745 47729 2773
rect 47763 2745 47791 2773
rect 47577 876 47605 904
rect 47639 876 47667 904
rect 47701 876 47729 904
rect 47763 876 47791 904
rect 47577 814 47605 842
rect 47639 814 47667 842
rect 47701 814 47729 842
rect 47763 814 47791 842
rect 47577 752 47605 780
rect 47639 752 47667 780
rect 47701 752 47729 780
rect 47763 752 47791 780
rect 47577 690 47605 718
rect 47639 690 47667 718
rect 47701 690 47729 718
rect 47763 690 47791 718
rect 49437 5931 49465 5959
rect 49499 5931 49527 5959
rect 49561 5931 49589 5959
rect 49623 5931 49651 5959
rect 49437 5869 49465 5897
rect 49499 5869 49527 5897
rect 49561 5869 49589 5897
rect 49623 5869 49651 5897
rect 49437 5807 49465 5835
rect 49499 5807 49527 5835
rect 49561 5807 49589 5835
rect 49623 5807 49651 5835
rect 49437 5745 49465 5773
rect 49499 5745 49527 5773
rect 49561 5745 49589 5773
rect 49623 5745 49651 5773
rect 49437 396 49465 424
rect 49499 396 49527 424
rect 49561 396 49589 424
rect 49623 396 49651 424
rect 49437 334 49465 362
rect 49499 334 49527 362
rect 49561 334 49589 362
rect 49623 334 49651 362
rect 49437 272 49465 300
rect 49499 272 49527 300
rect 49561 272 49589 300
rect 49623 272 49651 300
rect 49437 210 49465 238
rect 49499 210 49527 238
rect 49561 210 49589 238
rect 49623 210 49651 238
rect 56577 11931 56605 11959
rect 56639 11931 56667 11959
rect 56701 11931 56729 11959
rect 56763 11931 56791 11959
rect 56577 11869 56605 11897
rect 56639 11869 56667 11897
rect 56701 11869 56729 11897
rect 56763 11869 56791 11897
rect 56577 11807 56605 11835
rect 56639 11807 56667 11835
rect 56701 11807 56729 11835
rect 56763 11807 56791 11835
rect 56577 11745 56605 11773
rect 56639 11745 56667 11773
rect 56701 11745 56729 11773
rect 56763 11745 56791 11773
rect 56577 2931 56605 2959
rect 56639 2931 56667 2959
rect 56701 2931 56729 2959
rect 56763 2931 56791 2959
rect 56577 2869 56605 2897
rect 56639 2869 56667 2897
rect 56701 2869 56729 2897
rect 56763 2869 56791 2897
rect 56577 2807 56605 2835
rect 56639 2807 56667 2835
rect 56701 2807 56729 2835
rect 56763 2807 56791 2835
rect 56577 2745 56605 2773
rect 56639 2745 56667 2773
rect 56701 2745 56729 2773
rect 56763 2745 56791 2773
rect 56577 876 56605 904
rect 56639 876 56667 904
rect 56701 876 56729 904
rect 56763 876 56791 904
rect 56577 814 56605 842
rect 56639 814 56667 842
rect 56701 814 56729 842
rect 56763 814 56791 842
rect 56577 752 56605 780
rect 56639 752 56667 780
rect 56701 752 56729 780
rect 56763 752 56791 780
rect 56577 690 56605 718
rect 56639 690 56667 718
rect 56701 690 56729 718
rect 56763 690 56791 718
rect 58437 5931 58465 5959
rect 58499 5931 58527 5959
rect 58561 5931 58589 5959
rect 58623 5931 58651 5959
rect 58437 5869 58465 5897
rect 58499 5869 58527 5897
rect 58561 5869 58589 5897
rect 58623 5869 58651 5897
rect 58437 5807 58465 5835
rect 58499 5807 58527 5835
rect 58561 5807 58589 5835
rect 58623 5807 58651 5835
rect 58437 5745 58465 5773
rect 58499 5745 58527 5773
rect 58561 5745 58589 5773
rect 58623 5745 58651 5773
rect 58437 396 58465 424
rect 58499 396 58527 424
rect 58561 396 58589 424
rect 58623 396 58651 424
rect 58437 334 58465 362
rect 58499 334 58527 362
rect 58561 334 58589 362
rect 58623 334 58651 362
rect 58437 272 58465 300
rect 58499 272 58527 300
rect 58561 272 58589 300
rect 58623 272 58651 300
rect 58437 210 58465 238
rect 58499 210 58527 238
rect 58561 210 58589 238
rect 58623 210 58651 238
rect 65577 11931 65605 11959
rect 65639 11931 65667 11959
rect 65701 11931 65729 11959
rect 65763 11931 65791 11959
rect 65577 11869 65605 11897
rect 65639 11869 65667 11897
rect 65701 11869 65729 11897
rect 65763 11869 65791 11897
rect 65577 11807 65605 11835
rect 65639 11807 65667 11835
rect 65701 11807 65729 11835
rect 65763 11807 65791 11835
rect 65577 11745 65605 11773
rect 65639 11745 65667 11773
rect 65701 11745 65729 11773
rect 65763 11745 65791 11773
rect 65577 2931 65605 2959
rect 65639 2931 65667 2959
rect 65701 2931 65729 2959
rect 65763 2931 65791 2959
rect 65577 2869 65605 2897
rect 65639 2869 65667 2897
rect 65701 2869 65729 2897
rect 65763 2869 65791 2897
rect 65577 2807 65605 2835
rect 65639 2807 65667 2835
rect 65701 2807 65729 2835
rect 65763 2807 65791 2835
rect 65577 2745 65605 2773
rect 65639 2745 65667 2773
rect 65701 2745 65729 2773
rect 65763 2745 65791 2773
rect 65577 876 65605 904
rect 65639 876 65667 904
rect 65701 876 65729 904
rect 65763 876 65791 904
rect 65577 814 65605 842
rect 65639 814 65667 842
rect 65701 814 65729 842
rect 65763 814 65791 842
rect 65577 752 65605 780
rect 65639 752 65667 780
rect 65701 752 65729 780
rect 65763 752 65791 780
rect 65577 690 65605 718
rect 65639 690 65667 718
rect 65701 690 65729 718
rect 65763 690 65791 718
rect 67437 5931 67465 5959
rect 67499 5931 67527 5959
rect 67561 5931 67589 5959
rect 67623 5931 67651 5959
rect 67437 5869 67465 5897
rect 67499 5869 67527 5897
rect 67561 5869 67589 5897
rect 67623 5869 67651 5897
rect 67437 5807 67465 5835
rect 67499 5807 67527 5835
rect 67561 5807 67589 5835
rect 67623 5807 67651 5835
rect 67437 5745 67465 5773
rect 67499 5745 67527 5773
rect 67561 5745 67589 5773
rect 67623 5745 67651 5773
rect 67437 396 67465 424
rect 67499 396 67527 424
rect 67561 396 67589 424
rect 67623 396 67651 424
rect 67437 334 67465 362
rect 67499 334 67527 362
rect 67561 334 67589 362
rect 67623 334 67651 362
rect 67437 272 67465 300
rect 67499 272 67527 300
rect 67561 272 67589 300
rect 67623 272 67651 300
rect 67437 210 67465 238
rect 67499 210 67527 238
rect 67561 210 67589 238
rect 67623 210 67651 238
rect 74577 11931 74605 11959
rect 74639 11931 74667 11959
rect 74701 11931 74729 11959
rect 74763 11931 74791 11959
rect 74577 11869 74605 11897
rect 74639 11869 74667 11897
rect 74701 11869 74729 11897
rect 74763 11869 74791 11897
rect 74577 11807 74605 11835
rect 74639 11807 74667 11835
rect 74701 11807 74729 11835
rect 74763 11807 74791 11835
rect 74577 11745 74605 11773
rect 74639 11745 74667 11773
rect 74701 11745 74729 11773
rect 74763 11745 74791 11773
rect 74577 2931 74605 2959
rect 74639 2931 74667 2959
rect 74701 2931 74729 2959
rect 74763 2931 74791 2959
rect 74577 2869 74605 2897
rect 74639 2869 74667 2897
rect 74701 2869 74729 2897
rect 74763 2869 74791 2897
rect 74577 2807 74605 2835
rect 74639 2807 74667 2835
rect 74701 2807 74729 2835
rect 74763 2807 74791 2835
rect 74577 2745 74605 2773
rect 74639 2745 74667 2773
rect 74701 2745 74729 2773
rect 74763 2745 74791 2773
rect 74577 876 74605 904
rect 74639 876 74667 904
rect 74701 876 74729 904
rect 74763 876 74791 904
rect 74577 814 74605 842
rect 74639 814 74667 842
rect 74701 814 74729 842
rect 74763 814 74791 842
rect 74577 752 74605 780
rect 74639 752 74667 780
rect 74701 752 74729 780
rect 74763 752 74791 780
rect 74577 690 74605 718
rect 74639 690 74667 718
rect 74701 690 74729 718
rect 74763 690 74791 718
rect 76437 5931 76465 5959
rect 76499 5931 76527 5959
rect 76561 5931 76589 5959
rect 76623 5931 76651 5959
rect 76437 5869 76465 5897
rect 76499 5869 76527 5897
rect 76561 5869 76589 5897
rect 76623 5869 76651 5897
rect 76437 5807 76465 5835
rect 76499 5807 76527 5835
rect 76561 5807 76589 5835
rect 76623 5807 76651 5835
rect 76437 5745 76465 5773
rect 76499 5745 76527 5773
rect 76561 5745 76589 5773
rect 76623 5745 76651 5773
rect 76437 396 76465 424
rect 76499 396 76527 424
rect 76561 396 76589 424
rect 76623 396 76651 424
rect 76437 334 76465 362
rect 76499 334 76527 362
rect 76561 334 76589 362
rect 76623 334 76651 362
rect 76437 272 76465 300
rect 76499 272 76527 300
rect 76561 272 76589 300
rect 76623 272 76651 300
rect 76437 210 76465 238
rect 76499 210 76527 238
rect 76561 210 76589 238
rect 76623 210 76651 238
rect 83577 11931 83605 11959
rect 83639 11931 83667 11959
rect 83701 11931 83729 11959
rect 83763 11931 83791 11959
rect 83577 11869 83605 11897
rect 83639 11869 83667 11897
rect 83701 11869 83729 11897
rect 83763 11869 83791 11897
rect 83577 11807 83605 11835
rect 83639 11807 83667 11835
rect 83701 11807 83729 11835
rect 83763 11807 83791 11835
rect 83577 11745 83605 11773
rect 83639 11745 83667 11773
rect 83701 11745 83729 11773
rect 83763 11745 83791 11773
rect 83577 2931 83605 2959
rect 83639 2931 83667 2959
rect 83701 2931 83729 2959
rect 83763 2931 83791 2959
rect 83577 2869 83605 2897
rect 83639 2869 83667 2897
rect 83701 2869 83729 2897
rect 83763 2869 83791 2897
rect 83577 2807 83605 2835
rect 83639 2807 83667 2835
rect 83701 2807 83729 2835
rect 83763 2807 83791 2835
rect 83577 2745 83605 2773
rect 83639 2745 83667 2773
rect 83701 2745 83729 2773
rect 83763 2745 83791 2773
rect 83577 876 83605 904
rect 83639 876 83667 904
rect 83701 876 83729 904
rect 83763 876 83791 904
rect 83577 814 83605 842
rect 83639 814 83667 842
rect 83701 814 83729 842
rect 83763 814 83791 842
rect 83577 752 83605 780
rect 83639 752 83667 780
rect 83701 752 83729 780
rect 83763 752 83791 780
rect 83577 690 83605 718
rect 83639 690 83667 718
rect 83701 690 83729 718
rect 83763 690 83791 718
rect 85437 5931 85465 5959
rect 85499 5931 85527 5959
rect 85561 5931 85589 5959
rect 85623 5931 85651 5959
rect 85437 5869 85465 5897
rect 85499 5869 85527 5897
rect 85561 5869 85589 5897
rect 85623 5869 85651 5897
rect 85437 5807 85465 5835
rect 85499 5807 85527 5835
rect 85561 5807 85589 5835
rect 85623 5807 85651 5835
rect 85437 5745 85465 5773
rect 85499 5745 85527 5773
rect 85561 5745 85589 5773
rect 85623 5745 85651 5773
rect 85437 396 85465 424
rect 85499 396 85527 424
rect 85561 396 85589 424
rect 85623 396 85651 424
rect 85437 334 85465 362
rect 85499 334 85527 362
rect 85561 334 85589 362
rect 85623 334 85651 362
rect 85437 272 85465 300
rect 85499 272 85527 300
rect 85561 272 85589 300
rect 85623 272 85651 300
rect 85437 210 85465 238
rect 85499 210 85527 238
rect 85561 210 85589 238
rect 85623 210 85651 238
rect 92577 11931 92605 11959
rect 92639 11931 92667 11959
rect 92701 11931 92729 11959
rect 92763 11931 92791 11959
rect 92577 11869 92605 11897
rect 92639 11869 92667 11897
rect 92701 11869 92729 11897
rect 92763 11869 92791 11897
rect 92577 11807 92605 11835
rect 92639 11807 92667 11835
rect 92701 11807 92729 11835
rect 92763 11807 92791 11835
rect 92577 11745 92605 11773
rect 92639 11745 92667 11773
rect 92701 11745 92729 11773
rect 92763 11745 92791 11773
rect 92577 2931 92605 2959
rect 92639 2931 92667 2959
rect 92701 2931 92729 2959
rect 92763 2931 92791 2959
rect 92577 2869 92605 2897
rect 92639 2869 92667 2897
rect 92701 2869 92729 2897
rect 92763 2869 92791 2897
rect 92577 2807 92605 2835
rect 92639 2807 92667 2835
rect 92701 2807 92729 2835
rect 92763 2807 92791 2835
rect 92577 2745 92605 2773
rect 92639 2745 92667 2773
rect 92701 2745 92729 2773
rect 92763 2745 92791 2773
rect 92577 876 92605 904
rect 92639 876 92667 904
rect 92701 876 92729 904
rect 92763 876 92791 904
rect 92577 814 92605 842
rect 92639 814 92667 842
rect 92701 814 92729 842
rect 92763 814 92791 842
rect 92577 752 92605 780
rect 92639 752 92667 780
rect 92701 752 92729 780
rect 92763 752 92791 780
rect 92577 690 92605 718
rect 92639 690 92667 718
rect 92701 690 92729 718
rect 92763 690 92791 718
rect 94437 5931 94465 5959
rect 94499 5931 94527 5959
rect 94561 5931 94589 5959
rect 94623 5931 94651 5959
rect 94437 5869 94465 5897
rect 94499 5869 94527 5897
rect 94561 5869 94589 5897
rect 94623 5869 94651 5897
rect 94437 5807 94465 5835
rect 94499 5807 94527 5835
rect 94561 5807 94589 5835
rect 94623 5807 94651 5835
rect 94437 5745 94465 5773
rect 94499 5745 94527 5773
rect 94561 5745 94589 5773
rect 94623 5745 94651 5773
rect 94437 396 94465 424
rect 94499 396 94527 424
rect 94561 396 94589 424
rect 94623 396 94651 424
rect 94437 334 94465 362
rect 94499 334 94527 362
rect 94561 334 94589 362
rect 94623 334 94651 362
rect 94437 272 94465 300
rect 94499 272 94527 300
rect 94561 272 94589 300
rect 94623 272 94651 300
rect 94437 210 94465 238
rect 94499 210 94527 238
rect 94561 210 94589 238
rect 94623 210 94651 238
rect 101577 11931 101605 11959
rect 101639 11931 101667 11959
rect 101701 11931 101729 11959
rect 101763 11931 101791 11959
rect 101577 11869 101605 11897
rect 101639 11869 101667 11897
rect 101701 11869 101729 11897
rect 101763 11869 101791 11897
rect 101577 11807 101605 11835
rect 101639 11807 101667 11835
rect 101701 11807 101729 11835
rect 101763 11807 101791 11835
rect 101577 11745 101605 11773
rect 101639 11745 101667 11773
rect 101701 11745 101729 11773
rect 101763 11745 101791 11773
rect 101577 2931 101605 2959
rect 101639 2931 101667 2959
rect 101701 2931 101729 2959
rect 101763 2931 101791 2959
rect 101577 2869 101605 2897
rect 101639 2869 101667 2897
rect 101701 2869 101729 2897
rect 101763 2869 101791 2897
rect 101577 2807 101605 2835
rect 101639 2807 101667 2835
rect 101701 2807 101729 2835
rect 101763 2807 101791 2835
rect 101577 2745 101605 2773
rect 101639 2745 101667 2773
rect 101701 2745 101729 2773
rect 101763 2745 101791 2773
rect 101577 876 101605 904
rect 101639 876 101667 904
rect 101701 876 101729 904
rect 101763 876 101791 904
rect 101577 814 101605 842
rect 101639 814 101667 842
rect 101701 814 101729 842
rect 101763 814 101791 842
rect 101577 752 101605 780
rect 101639 752 101667 780
rect 101701 752 101729 780
rect 101763 752 101791 780
rect 101577 690 101605 718
rect 101639 690 101667 718
rect 101701 690 101729 718
rect 101763 690 101791 718
rect 103437 5931 103465 5959
rect 103499 5931 103527 5959
rect 103561 5931 103589 5959
rect 103623 5931 103651 5959
rect 103437 5869 103465 5897
rect 103499 5869 103527 5897
rect 103561 5869 103589 5897
rect 103623 5869 103651 5897
rect 103437 5807 103465 5835
rect 103499 5807 103527 5835
rect 103561 5807 103589 5835
rect 103623 5807 103651 5835
rect 103437 5745 103465 5773
rect 103499 5745 103527 5773
rect 103561 5745 103589 5773
rect 103623 5745 103651 5773
rect 103437 396 103465 424
rect 103499 396 103527 424
rect 103561 396 103589 424
rect 103623 396 103651 424
rect 103437 334 103465 362
rect 103499 334 103527 362
rect 103561 334 103589 362
rect 103623 334 103651 362
rect 103437 272 103465 300
rect 103499 272 103527 300
rect 103561 272 103589 300
rect 103623 272 103651 300
rect 103437 210 103465 238
rect 103499 210 103527 238
rect 103561 210 103589 238
rect 103623 210 103651 238
rect 110577 11931 110605 11959
rect 110639 11931 110667 11959
rect 110701 11931 110729 11959
rect 110763 11931 110791 11959
rect 110577 11869 110605 11897
rect 110639 11869 110667 11897
rect 110701 11869 110729 11897
rect 110763 11869 110791 11897
rect 110577 11807 110605 11835
rect 110639 11807 110667 11835
rect 110701 11807 110729 11835
rect 110763 11807 110791 11835
rect 110577 11745 110605 11773
rect 110639 11745 110667 11773
rect 110701 11745 110729 11773
rect 110763 11745 110791 11773
rect 110577 2931 110605 2959
rect 110639 2931 110667 2959
rect 110701 2931 110729 2959
rect 110763 2931 110791 2959
rect 110577 2869 110605 2897
rect 110639 2869 110667 2897
rect 110701 2869 110729 2897
rect 110763 2869 110791 2897
rect 110577 2807 110605 2835
rect 110639 2807 110667 2835
rect 110701 2807 110729 2835
rect 110763 2807 110791 2835
rect 110577 2745 110605 2773
rect 110639 2745 110667 2773
rect 110701 2745 110729 2773
rect 110763 2745 110791 2773
rect 110577 876 110605 904
rect 110639 876 110667 904
rect 110701 876 110729 904
rect 110763 876 110791 904
rect 110577 814 110605 842
rect 110639 814 110667 842
rect 110701 814 110729 842
rect 110763 814 110791 842
rect 110577 752 110605 780
rect 110639 752 110667 780
rect 110701 752 110729 780
rect 110763 752 110791 780
rect 110577 690 110605 718
rect 110639 690 110667 718
rect 110701 690 110729 718
rect 110763 690 110791 718
rect 112437 5931 112465 5959
rect 112499 5931 112527 5959
rect 112561 5931 112589 5959
rect 112623 5931 112651 5959
rect 112437 5869 112465 5897
rect 112499 5869 112527 5897
rect 112561 5869 112589 5897
rect 112623 5869 112651 5897
rect 112437 5807 112465 5835
rect 112499 5807 112527 5835
rect 112561 5807 112589 5835
rect 112623 5807 112651 5835
rect 112437 5745 112465 5773
rect 112499 5745 112527 5773
rect 112561 5745 112589 5773
rect 112623 5745 112651 5773
rect 112437 396 112465 424
rect 112499 396 112527 424
rect 112561 396 112589 424
rect 112623 396 112651 424
rect 112437 334 112465 362
rect 112499 334 112527 362
rect 112561 334 112589 362
rect 112623 334 112651 362
rect 112437 272 112465 300
rect 112499 272 112527 300
rect 112561 272 112589 300
rect 112623 272 112651 300
rect 112437 210 112465 238
rect 112499 210 112527 238
rect 112561 210 112589 238
rect 112623 210 112651 238
rect 119577 11931 119605 11959
rect 119639 11931 119667 11959
rect 119701 11931 119729 11959
rect 119763 11931 119791 11959
rect 119577 11869 119605 11897
rect 119639 11869 119667 11897
rect 119701 11869 119729 11897
rect 119763 11869 119791 11897
rect 119577 11807 119605 11835
rect 119639 11807 119667 11835
rect 119701 11807 119729 11835
rect 119763 11807 119791 11835
rect 119577 11745 119605 11773
rect 119639 11745 119667 11773
rect 119701 11745 119729 11773
rect 119763 11745 119791 11773
rect 119577 2931 119605 2959
rect 119639 2931 119667 2959
rect 119701 2931 119729 2959
rect 119763 2931 119791 2959
rect 119577 2869 119605 2897
rect 119639 2869 119667 2897
rect 119701 2869 119729 2897
rect 119763 2869 119791 2897
rect 119577 2807 119605 2835
rect 119639 2807 119667 2835
rect 119701 2807 119729 2835
rect 119763 2807 119791 2835
rect 119577 2745 119605 2773
rect 119639 2745 119667 2773
rect 119701 2745 119729 2773
rect 119763 2745 119791 2773
rect 119577 876 119605 904
rect 119639 876 119667 904
rect 119701 876 119729 904
rect 119763 876 119791 904
rect 119577 814 119605 842
rect 119639 814 119667 842
rect 119701 814 119729 842
rect 119763 814 119791 842
rect 119577 752 119605 780
rect 119639 752 119667 780
rect 119701 752 119729 780
rect 119763 752 119791 780
rect 119577 690 119605 718
rect 119639 690 119667 718
rect 119701 690 119729 718
rect 119763 690 119791 718
rect 121437 5931 121465 5959
rect 121499 5931 121527 5959
rect 121561 5931 121589 5959
rect 121623 5931 121651 5959
rect 121437 5869 121465 5897
rect 121499 5869 121527 5897
rect 121561 5869 121589 5897
rect 121623 5869 121651 5897
rect 121437 5807 121465 5835
rect 121499 5807 121527 5835
rect 121561 5807 121589 5835
rect 121623 5807 121651 5835
rect 121437 5745 121465 5773
rect 121499 5745 121527 5773
rect 121561 5745 121589 5773
rect 121623 5745 121651 5773
rect 121437 396 121465 424
rect 121499 396 121527 424
rect 121561 396 121589 424
rect 121623 396 121651 424
rect 121437 334 121465 362
rect 121499 334 121527 362
rect 121561 334 121589 362
rect 121623 334 121651 362
rect 121437 272 121465 300
rect 121499 272 121527 300
rect 121561 272 121589 300
rect 121623 272 121651 300
rect 121437 210 121465 238
rect 121499 210 121527 238
rect 121561 210 121589 238
rect 121623 210 121651 238
rect 128577 11931 128605 11959
rect 128639 11931 128667 11959
rect 128701 11931 128729 11959
rect 128763 11931 128791 11959
rect 128577 11869 128605 11897
rect 128639 11869 128667 11897
rect 128701 11869 128729 11897
rect 128763 11869 128791 11897
rect 128577 11807 128605 11835
rect 128639 11807 128667 11835
rect 128701 11807 128729 11835
rect 128763 11807 128791 11835
rect 128577 11745 128605 11773
rect 128639 11745 128667 11773
rect 128701 11745 128729 11773
rect 128763 11745 128791 11773
rect 128577 2931 128605 2959
rect 128639 2931 128667 2959
rect 128701 2931 128729 2959
rect 128763 2931 128791 2959
rect 128577 2869 128605 2897
rect 128639 2869 128667 2897
rect 128701 2869 128729 2897
rect 128763 2869 128791 2897
rect 128577 2807 128605 2835
rect 128639 2807 128667 2835
rect 128701 2807 128729 2835
rect 128763 2807 128791 2835
rect 128577 2745 128605 2773
rect 128639 2745 128667 2773
rect 128701 2745 128729 2773
rect 128763 2745 128791 2773
rect 128577 876 128605 904
rect 128639 876 128667 904
rect 128701 876 128729 904
rect 128763 876 128791 904
rect 128577 814 128605 842
rect 128639 814 128667 842
rect 128701 814 128729 842
rect 128763 814 128791 842
rect 128577 752 128605 780
rect 128639 752 128667 780
rect 128701 752 128729 780
rect 128763 752 128791 780
rect 128577 690 128605 718
rect 128639 690 128667 718
rect 128701 690 128729 718
rect 128763 690 128791 718
rect 130437 5931 130465 5959
rect 130499 5931 130527 5959
rect 130561 5931 130589 5959
rect 130623 5931 130651 5959
rect 130437 5869 130465 5897
rect 130499 5869 130527 5897
rect 130561 5869 130589 5897
rect 130623 5869 130651 5897
rect 130437 5807 130465 5835
rect 130499 5807 130527 5835
rect 130561 5807 130589 5835
rect 130623 5807 130651 5835
rect 130437 5745 130465 5773
rect 130499 5745 130527 5773
rect 130561 5745 130589 5773
rect 130623 5745 130651 5773
rect 130437 396 130465 424
rect 130499 396 130527 424
rect 130561 396 130589 424
rect 130623 396 130651 424
rect 130437 334 130465 362
rect 130499 334 130527 362
rect 130561 334 130589 362
rect 130623 334 130651 362
rect 130437 272 130465 300
rect 130499 272 130527 300
rect 130561 272 130589 300
rect 130623 272 130651 300
rect 130437 210 130465 238
rect 130499 210 130527 238
rect 130561 210 130589 238
rect 130623 210 130651 238
rect 137577 11931 137605 11959
rect 137639 11931 137667 11959
rect 137701 11931 137729 11959
rect 137763 11931 137791 11959
rect 137577 11869 137605 11897
rect 137639 11869 137667 11897
rect 137701 11869 137729 11897
rect 137763 11869 137791 11897
rect 137577 11807 137605 11835
rect 137639 11807 137667 11835
rect 137701 11807 137729 11835
rect 137763 11807 137791 11835
rect 137577 11745 137605 11773
rect 137639 11745 137667 11773
rect 137701 11745 137729 11773
rect 137763 11745 137791 11773
rect 137577 2931 137605 2959
rect 137639 2931 137667 2959
rect 137701 2931 137729 2959
rect 137763 2931 137791 2959
rect 137577 2869 137605 2897
rect 137639 2869 137667 2897
rect 137701 2869 137729 2897
rect 137763 2869 137791 2897
rect 137577 2807 137605 2835
rect 137639 2807 137667 2835
rect 137701 2807 137729 2835
rect 137763 2807 137791 2835
rect 137577 2745 137605 2773
rect 137639 2745 137667 2773
rect 137701 2745 137729 2773
rect 137763 2745 137791 2773
rect 137577 876 137605 904
rect 137639 876 137667 904
rect 137701 876 137729 904
rect 137763 876 137791 904
rect 137577 814 137605 842
rect 137639 814 137667 842
rect 137701 814 137729 842
rect 137763 814 137791 842
rect 137577 752 137605 780
rect 137639 752 137667 780
rect 137701 752 137729 780
rect 137763 752 137791 780
rect 137577 690 137605 718
rect 137639 690 137667 718
rect 137701 690 137729 718
rect 137763 690 137791 718
rect 139437 5931 139465 5959
rect 139499 5931 139527 5959
rect 139561 5931 139589 5959
rect 139623 5931 139651 5959
rect 139437 5869 139465 5897
rect 139499 5869 139527 5897
rect 139561 5869 139589 5897
rect 139623 5869 139651 5897
rect 139437 5807 139465 5835
rect 139499 5807 139527 5835
rect 139561 5807 139589 5835
rect 139623 5807 139651 5835
rect 139437 5745 139465 5773
rect 139499 5745 139527 5773
rect 139561 5745 139589 5773
rect 139623 5745 139651 5773
rect 139437 396 139465 424
rect 139499 396 139527 424
rect 139561 396 139589 424
rect 139623 396 139651 424
rect 139437 334 139465 362
rect 139499 334 139527 362
rect 139561 334 139589 362
rect 139623 334 139651 362
rect 139437 272 139465 300
rect 139499 272 139527 300
rect 139561 272 139589 300
rect 139623 272 139651 300
rect 139437 210 139465 238
rect 139499 210 139527 238
rect 139561 210 139589 238
rect 139623 210 139651 238
rect 146577 11931 146605 11959
rect 146639 11931 146667 11959
rect 146701 11931 146729 11959
rect 146763 11931 146791 11959
rect 146577 11869 146605 11897
rect 146639 11869 146667 11897
rect 146701 11869 146729 11897
rect 146763 11869 146791 11897
rect 146577 11807 146605 11835
rect 146639 11807 146667 11835
rect 146701 11807 146729 11835
rect 146763 11807 146791 11835
rect 146577 11745 146605 11773
rect 146639 11745 146667 11773
rect 146701 11745 146729 11773
rect 146763 11745 146791 11773
rect 146577 2931 146605 2959
rect 146639 2931 146667 2959
rect 146701 2931 146729 2959
rect 146763 2931 146791 2959
rect 146577 2869 146605 2897
rect 146639 2869 146667 2897
rect 146701 2869 146729 2897
rect 146763 2869 146791 2897
rect 146577 2807 146605 2835
rect 146639 2807 146667 2835
rect 146701 2807 146729 2835
rect 146763 2807 146791 2835
rect 146577 2745 146605 2773
rect 146639 2745 146667 2773
rect 146701 2745 146729 2773
rect 146763 2745 146791 2773
rect 146577 876 146605 904
rect 146639 876 146667 904
rect 146701 876 146729 904
rect 146763 876 146791 904
rect 146577 814 146605 842
rect 146639 814 146667 842
rect 146701 814 146729 842
rect 146763 814 146791 842
rect 146577 752 146605 780
rect 146639 752 146667 780
rect 146701 752 146729 780
rect 146763 752 146791 780
rect 146577 690 146605 718
rect 146639 690 146667 718
rect 146701 690 146729 718
rect 146763 690 146791 718
rect 148437 5931 148465 5959
rect 148499 5931 148527 5959
rect 148561 5931 148589 5959
rect 148623 5931 148651 5959
rect 148437 5869 148465 5897
rect 148499 5869 148527 5897
rect 148561 5869 148589 5897
rect 148623 5869 148651 5897
rect 148437 5807 148465 5835
rect 148499 5807 148527 5835
rect 148561 5807 148589 5835
rect 148623 5807 148651 5835
rect 148437 5745 148465 5773
rect 148499 5745 148527 5773
rect 148561 5745 148589 5773
rect 148623 5745 148651 5773
rect 148437 396 148465 424
rect 148499 396 148527 424
rect 148561 396 148589 424
rect 148623 396 148651 424
rect 148437 334 148465 362
rect 148499 334 148527 362
rect 148561 334 148589 362
rect 148623 334 148651 362
rect 148437 272 148465 300
rect 148499 272 148527 300
rect 148561 272 148589 300
rect 148623 272 148651 300
rect 148437 210 148465 238
rect 148499 210 148527 238
rect 148561 210 148589 238
rect 148623 210 148651 238
rect 155577 11931 155605 11959
rect 155639 11931 155667 11959
rect 155701 11931 155729 11959
rect 155763 11931 155791 11959
rect 155577 11869 155605 11897
rect 155639 11869 155667 11897
rect 155701 11869 155729 11897
rect 155763 11869 155791 11897
rect 155577 11807 155605 11835
rect 155639 11807 155667 11835
rect 155701 11807 155729 11835
rect 155763 11807 155791 11835
rect 155577 11745 155605 11773
rect 155639 11745 155667 11773
rect 155701 11745 155729 11773
rect 155763 11745 155791 11773
rect 155577 2931 155605 2959
rect 155639 2931 155667 2959
rect 155701 2931 155729 2959
rect 155763 2931 155791 2959
rect 155577 2869 155605 2897
rect 155639 2869 155667 2897
rect 155701 2869 155729 2897
rect 155763 2869 155791 2897
rect 155577 2807 155605 2835
rect 155639 2807 155667 2835
rect 155701 2807 155729 2835
rect 155763 2807 155791 2835
rect 155577 2745 155605 2773
rect 155639 2745 155667 2773
rect 155701 2745 155729 2773
rect 155763 2745 155791 2773
rect 155577 876 155605 904
rect 155639 876 155667 904
rect 155701 876 155729 904
rect 155763 876 155791 904
rect 155577 814 155605 842
rect 155639 814 155667 842
rect 155701 814 155729 842
rect 155763 814 155791 842
rect 155577 752 155605 780
rect 155639 752 155667 780
rect 155701 752 155729 780
rect 155763 752 155791 780
rect 155577 690 155605 718
rect 155639 690 155667 718
rect 155701 690 155729 718
rect 155763 690 155791 718
rect 157437 5931 157465 5959
rect 157499 5931 157527 5959
rect 157561 5931 157589 5959
rect 157623 5931 157651 5959
rect 157437 5869 157465 5897
rect 157499 5869 157527 5897
rect 157561 5869 157589 5897
rect 157623 5869 157651 5897
rect 157437 5807 157465 5835
rect 157499 5807 157527 5835
rect 157561 5807 157589 5835
rect 157623 5807 157651 5835
rect 157437 5745 157465 5773
rect 157499 5745 157527 5773
rect 157561 5745 157589 5773
rect 157623 5745 157651 5773
rect 157437 396 157465 424
rect 157499 396 157527 424
rect 157561 396 157589 424
rect 157623 396 157651 424
rect 157437 334 157465 362
rect 157499 334 157527 362
rect 157561 334 157589 362
rect 157623 334 157651 362
rect 157437 272 157465 300
rect 157499 272 157527 300
rect 157561 272 157589 300
rect 157623 272 157651 300
rect 157437 210 157465 238
rect 157499 210 157527 238
rect 157561 210 157589 238
rect 157623 210 157651 238
rect 164577 11931 164605 11959
rect 164639 11931 164667 11959
rect 164701 11931 164729 11959
rect 164763 11931 164791 11959
rect 164577 11869 164605 11897
rect 164639 11869 164667 11897
rect 164701 11869 164729 11897
rect 164763 11869 164791 11897
rect 164577 11807 164605 11835
rect 164639 11807 164667 11835
rect 164701 11807 164729 11835
rect 164763 11807 164791 11835
rect 164577 11745 164605 11773
rect 164639 11745 164667 11773
rect 164701 11745 164729 11773
rect 164763 11745 164791 11773
rect 164577 2931 164605 2959
rect 164639 2931 164667 2959
rect 164701 2931 164729 2959
rect 164763 2931 164791 2959
rect 164577 2869 164605 2897
rect 164639 2869 164667 2897
rect 164701 2869 164729 2897
rect 164763 2869 164791 2897
rect 164577 2807 164605 2835
rect 164639 2807 164667 2835
rect 164701 2807 164729 2835
rect 164763 2807 164791 2835
rect 164577 2745 164605 2773
rect 164639 2745 164667 2773
rect 164701 2745 164729 2773
rect 164763 2745 164791 2773
rect 164577 876 164605 904
rect 164639 876 164667 904
rect 164701 876 164729 904
rect 164763 876 164791 904
rect 164577 814 164605 842
rect 164639 814 164667 842
rect 164701 814 164729 842
rect 164763 814 164791 842
rect 164577 752 164605 780
rect 164639 752 164667 780
rect 164701 752 164729 780
rect 164763 752 164791 780
rect 164577 690 164605 718
rect 164639 690 164667 718
rect 164701 690 164729 718
rect 164763 690 164791 718
rect 166437 5931 166465 5959
rect 166499 5931 166527 5959
rect 166561 5931 166589 5959
rect 166623 5931 166651 5959
rect 166437 5869 166465 5897
rect 166499 5869 166527 5897
rect 166561 5869 166589 5897
rect 166623 5869 166651 5897
rect 166437 5807 166465 5835
rect 166499 5807 166527 5835
rect 166561 5807 166589 5835
rect 166623 5807 166651 5835
rect 166437 5745 166465 5773
rect 166499 5745 166527 5773
rect 166561 5745 166589 5773
rect 166623 5745 166651 5773
rect 166437 396 166465 424
rect 166499 396 166527 424
rect 166561 396 166589 424
rect 166623 396 166651 424
rect 166437 334 166465 362
rect 166499 334 166527 362
rect 166561 334 166589 362
rect 166623 334 166651 362
rect 166437 272 166465 300
rect 166499 272 166527 300
rect 166561 272 166589 300
rect 166623 272 166651 300
rect 166437 210 166465 238
rect 166499 210 166527 238
rect 166561 210 166589 238
rect 166623 210 166651 238
rect 173577 11931 173605 11959
rect 173639 11931 173667 11959
rect 173701 11931 173729 11959
rect 173763 11931 173791 11959
rect 173577 11869 173605 11897
rect 173639 11869 173667 11897
rect 173701 11869 173729 11897
rect 173763 11869 173791 11897
rect 173577 11807 173605 11835
rect 173639 11807 173667 11835
rect 173701 11807 173729 11835
rect 173763 11807 173791 11835
rect 173577 11745 173605 11773
rect 173639 11745 173667 11773
rect 173701 11745 173729 11773
rect 173763 11745 173791 11773
rect 173577 2931 173605 2959
rect 173639 2931 173667 2959
rect 173701 2931 173729 2959
rect 173763 2931 173791 2959
rect 173577 2869 173605 2897
rect 173639 2869 173667 2897
rect 173701 2869 173729 2897
rect 173763 2869 173791 2897
rect 173577 2807 173605 2835
rect 173639 2807 173667 2835
rect 173701 2807 173729 2835
rect 173763 2807 173791 2835
rect 173577 2745 173605 2773
rect 173639 2745 173667 2773
rect 173701 2745 173729 2773
rect 173763 2745 173791 2773
rect 173577 876 173605 904
rect 173639 876 173667 904
rect 173701 876 173729 904
rect 173763 876 173791 904
rect 173577 814 173605 842
rect 173639 814 173667 842
rect 173701 814 173729 842
rect 173763 814 173791 842
rect 173577 752 173605 780
rect 173639 752 173667 780
rect 173701 752 173729 780
rect 173763 752 173791 780
rect 173577 690 173605 718
rect 173639 690 173667 718
rect 173701 690 173729 718
rect 173763 690 173791 718
rect 175437 5931 175465 5959
rect 175499 5931 175527 5959
rect 175561 5931 175589 5959
rect 175623 5931 175651 5959
rect 175437 5869 175465 5897
rect 175499 5869 175527 5897
rect 175561 5869 175589 5897
rect 175623 5869 175651 5897
rect 175437 5807 175465 5835
rect 175499 5807 175527 5835
rect 175561 5807 175589 5835
rect 175623 5807 175651 5835
rect 175437 5745 175465 5773
rect 175499 5745 175527 5773
rect 175561 5745 175589 5773
rect 175623 5745 175651 5773
rect 175437 396 175465 424
rect 175499 396 175527 424
rect 175561 396 175589 424
rect 175623 396 175651 424
rect 175437 334 175465 362
rect 175499 334 175527 362
rect 175561 334 175589 362
rect 175623 334 175651 362
rect 175437 272 175465 300
rect 175499 272 175527 300
rect 175561 272 175589 300
rect 175623 272 175651 300
rect 175437 210 175465 238
rect 175499 210 175527 238
rect 175561 210 175589 238
rect 175623 210 175651 238
rect 182577 11931 182605 11959
rect 182639 11931 182667 11959
rect 182701 11931 182729 11959
rect 182763 11931 182791 11959
rect 182577 11869 182605 11897
rect 182639 11869 182667 11897
rect 182701 11869 182729 11897
rect 182763 11869 182791 11897
rect 182577 11807 182605 11835
rect 182639 11807 182667 11835
rect 182701 11807 182729 11835
rect 182763 11807 182791 11835
rect 182577 11745 182605 11773
rect 182639 11745 182667 11773
rect 182701 11745 182729 11773
rect 182763 11745 182791 11773
rect 182577 2931 182605 2959
rect 182639 2931 182667 2959
rect 182701 2931 182729 2959
rect 182763 2931 182791 2959
rect 182577 2869 182605 2897
rect 182639 2869 182667 2897
rect 182701 2869 182729 2897
rect 182763 2869 182791 2897
rect 182577 2807 182605 2835
rect 182639 2807 182667 2835
rect 182701 2807 182729 2835
rect 182763 2807 182791 2835
rect 182577 2745 182605 2773
rect 182639 2745 182667 2773
rect 182701 2745 182729 2773
rect 182763 2745 182791 2773
rect 182577 876 182605 904
rect 182639 876 182667 904
rect 182701 876 182729 904
rect 182763 876 182791 904
rect 182577 814 182605 842
rect 182639 814 182667 842
rect 182701 814 182729 842
rect 182763 814 182791 842
rect 182577 752 182605 780
rect 182639 752 182667 780
rect 182701 752 182729 780
rect 182763 752 182791 780
rect 182577 690 182605 718
rect 182639 690 182667 718
rect 182701 690 182729 718
rect 182763 690 182791 718
rect 184437 5931 184465 5959
rect 184499 5931 184527 5959
rect 184561 5931 184589 5959
rect 184623 5931 184651 5959
rect 184437 5869 184465 5897
rect 184499 5869 184527 5897
rect 184561 5869 184589 5897
rect 184623 5869 184651 5897
rect 184437 5807 184465 5835
rect 184499 5807 184527 5835
rect 184561 5807 184589 5835
rect 184623 5807 184651 5835
rect 184437 5745 184465 5773
rect 184499 5745 184527 5773
rect 184561 5745 184589 5773
rect 184623 5745 184651 5773
rect 184437 396 184465 424
rect 184499 396 184527 424
rect 184561 396 184589 424
rect 184623 396 184651 424
rect 184437 334 184465 362
rect 184499 334 184527 362
rect 184561 334 184589 362
rect 184623 334 184651 362
rect 184437 272 184465 300
rect 184499 272 184527 300
rect 184561 272 184589 300
rect 184623 272 184651 300
rect 184437 210 184465 238
rect 184499 210 184527 238
rect 184561 210 184589 238
rect 184623 210 184651 238
rect 191577 11931 191605 11959
rect 191639 11931 191667 11959
rect 191701 11931 191729 11959
rect 191763 11931 191791 11959
rect 191577 11869 191605 11897
rect 191639 11869 191667 11897
rect 191701 11869 191729 11897
rect 191763 11869 191791 11897
rect 191577 11807 191605 11835
rect 191639 11807 191667 11835
rect 191701 11807 191729 11835
rect 191763 11807 191791 11835
rect 191577 11745 191605 11773
rect 191639 11745 191667 11773
rect 191701 11745 191729 11773
rect 191763 11745 191791 11773
rect 191577 2931 191605 2959
rect 191639 2931 191667 2959
rect 191701 2931 191729 2959
rect 191763 2931 191791 2959
rect 191577 2869 191605 2897
rect 191639 2869 191667 2897
rect 191701 2869 191729 2897
rect 191763 2869 191791 2897
rect 191577 2807 191605 2835
rect 191639 2807 191667 2835
rect 191701 2807 191729 2835
rect 191763 2807 191791 2835
rect 191577 2745 191605 2773
rect 191639 2745 191667 2773
rect 191701 2745 191729 2773
rect 191763 2745 191791 2773
rect 191577 876 191605 904
rect 191639 876 191667 904
rect 191701 876 191729 904
rect 191763 876 191791 904
rect 191577 814 191605 842
rect 191639 814 191667 842
rect 191701 814 191729 842
rect 191763 814 191791 842
rect 191577 752 191605 780
rect 191639 752 191667 780
rect 191701 752 191729 780
rect 191763 752 191791 780
rect 191577 690 191605 718
rect 191639 690 191667 718
rect 191701 690 191729 718
rect 191763 690 191791 718
rect 193437 5931 193465 5959
rect 193499 5931 193527 5959
rect 193561 5931 193589 5959
rect 193623 5931 193651 5959
rect 193437 5869 193465 5897
rect 193499 5869 193527 5897
rect 193561 5869 193589 5897
rect 193623 5869 193651 5897
rect 193437 5807 193465 5835
rect 193499 5807 193527 5835
rect 193561 5807 193589 5835
rect 193623 5807 193651 5835
rect 193437 5745 193465 5773
rect 193499 5745 193527 5773
rect 193561 5745 193589 5773
rect 193623 5745 193651 5773
rect 193437 396 193465 424
rect 193499 396 193527 424
rect 193561 396 193589 424
rect 193623 396 193651 424
rect 193437 334 193465 362
rect 193499 334 193527 362
rect 193561 334 193589 362
rect 193623 334 193651 362
rect 193437 272 193465 300
rect 193499 272 193527 300
rect 193561 272 193589 300
rect 193623 272 193651 300
rect 193437 210 193465 238
rect 193499 210 193527 238
rect 193561 210 193589 238
rect 193623 210 193651 238
rect 200577 11931 200605 11959
rect 200639 11931 200667 11959
rect 200701 11931 200729 11959
rect 200763 11931 200791 11959
rect 200577 11869 200605 11897
rect 200639 11869 200667 11897
rect 200701 11869 200729 11897
rect 200763 11869 200791 11897
rect 200577 11807 200605 11835
rect 200639 11807 200667 11835
rect 200701 11807 200729 11835
rect 200763 11807 200791 11835
rect 200577 11745 200605 11773
rect 200639 11745 200667 11773
rect 200701 11745 200729 11773
rect 200763 11745 200791 11773
rect 200577 2931 200605 2959
rect 200639 2931 200667 2959
rect 200701 2931 200729 2959
rect 200763 2931 200791 2959
rect 200577 2869 200605 2897
rect 200639 2869 200667 2897
rect 200701 2869 200729 2897
rect 200763 2869 200791 2897
rect 200577 2807 200605 2835
rect 200639 2807 200667 2835
rect 200701 2807 200729 2835
rect 200763 2807 200791 2835
rect 200577 2745 200605 2773
rect 200639 2745 200667 2773
rect 200701 2745 200729 2773
rect 200763 2745 200791 2773
rect 200577 876 200605 904
rect 200639 876 200667 904
rect 200701 876 200729 904
rect 200763 876 200791 904
rect 200577 814 200605 842
rect 200639 814 200667 842
rect 200701 814 200729 842
rect 200763 814 200791 842
rect 200577 752 200605 780
rect 200639 752 200667 780
rect 200701 752 200729 780
rect 200763 752 200791 780
rect 200577 690 200605 718
rect 200639 690 200667 718
rect 200701 690 200729 718
rect 200763 690 200791 718
rect 202437 5931 202465 5959
rect 202499 5931 202527 5959
rect 202561 5931 202589 5959
rect 202623 5931 202651 5959
rect 202437 5869 202465 5897
rect 202499 5869 202527 5897
rect 202561 5869 202589 5897
rect 202623 5869 202651 5897
rect 202437 5807 202465 5835
rect 202499 5807 202527 5835
rect 202561 5807 202589 5835
rect 202623 5807 202651 5835
rect 202437 5745 202465 5773
rect 202499 5745 202527 5773
rect 202561 5745 202589 5773
rect 202623 5745 202651 5773
rect 202437 396 202465 424
rect 202499 396 202527 424
rect 202561 396 202589 424
rect 202623 396 202651 424
rect 202437 334 202465 362
rect 202499 334 202527 362
rect 202561 334 202589 362
rect 202623 334 202651 362
rect 202437 272 202465 300
rect 202499 272 202527 300
rect 202561 272 202589 300
rect 202623 272 202651 300
rect 202437 210 202465 238
rect 202499 210 202527 238
rect 202561 210 202589 238
rect 202623 210 202651 238
rect 209577 11931 209605 11959
rect 209639 11931 209667 11959
rect 209701 11931 209729 11959
rect 209763 11931 209791 11959
rect 209577 11869 209605 11897
rect 209639 11869 209667 11897
rect 209701 11869 209729 11897
rect 209763 11869 209791 11897
rect 209577 11807 209605 11835
rect 209639 11807 209667 11835
rect 209701 11807 209729 11835
rect 209763 11807 209791 11835
rect 209577 11745 209605 11773
rect 209639 11745 209667 11773
rect 209701 11745 209729 11773
rect 209763 11745 209791 11773
rect 209577 2931 209605 2959
rect 209639 2931 209667 2959
rect 209701 2931 209729 2959
rect 209763 2931 209791 2959
rect 209577 2869 209605 2897
rect 209639 2869 209667 2897
rect 209701 2869 209729 2897
rect 209763 2869 209791 2897
rect 209577 2807 209605 2835
rect 209639 2807 209667 2835
rect 209701 2807 209729 2835
rect 209763 2807 209791 2835
rect 209577 2745 209605 2773
rect 209639 2745 209667 2773
rect 209701 2745 209729 2773
rect 209763 2745 209791 2773
rect 209577 876 209605 904
rect 209639 876 209667 904
rect 209701 876 209729 904
rect 209763 876 209791 904
rect 209577 814 209605 842
rect 209639 814 209667 842
rect 209701 814 209729 842
rect 209763 814 209791 842
rect 209577 752 209605 780
rect 209639 752 209667 780
rect 209701 752 209729 780
rect 209763 752 209791 780
rect 209577 690 209605 718
rect 209639 690 209667 718
rect 209701 690 209729 718
rect 209763 690 209791 718
rect 211437 5931 211465 5959
rect 211499 5931 211527 5959
rect 211561 5931 211589 5959
rect 211623 5931 211651 5959
rect 211437 5869 211465 5897
rect 211499 5869 211527 5897
rect 211561 5869 211589 5897
rect 211623 5869 211651 5897
rect 211437 5807 211465 5835
rect 211499 5807 211527 5835
rect 211561 5807 211589 5835
rect 211623 5807 211651 5835
rect 211437 5745 211465 5773
rect 211499 5745 211527 5773
rect 211561 5745 211589 5773
rect 211623 5745 211651 5773
rect 211437 396 211465 424
rect 211499 396 211527 424
rect 211561 396 211589 424
rect 211623 396 211651 424
rect 211437 334 211465 362
rect 211499 334 211527 362
rect 211561 334 211589 362
rect 211623 334 211651 362
rect 211437 272 211465 300
rect 211499 272 211527 300
rect 211561 272 211589 300
rect 211623 272 211651 300
rect 211437 210 211465 238
rect 211499 210 211527 238
rect 211561 210 211589 238
rect 211623 210 211651 238
rect 218577 11931 218605 11959
rect 218639 11931 218667 11959
rect 218701 11931 218729 11959
rect 218763 11931 218791 11959
rect 218577 11869 218605 11897
rect 218639 11869 218667 11897
rect 218701 11869 218729 11897
rect 218763 11869 218791 11897
rect 218577 11807 218605 11835
rect 218639 11807 218667 11835
rect 218701 11807 218729 11835
rect 218763 11807 218791 11835
rect 218577 11745 218605 11773
rect 218639 11745 218667 11773
rect 218701 11745 218729 11773
rect 218763 11745 218791 11773
rect 218577 2931 218605 2959
rect 218639 2931 218667 2959
rect 218701 2931 218729 2959
rect 218763 2931 218791 2959
rect 218577 2869 218605 2897
rect 218639 2869 218667 2897
rect 218701 2869 218729 2897
rect 218763 2869 218791 2897
rect 218577 2807 218605 2835
rect 218639 2807 218667 2835
rect 218701 2807 218729 2835
rect 218763 2807 218791 2835
rect 218577 2745 218605 2773
rect 218639 2745 218667 2773
rect 218701 2745 218729 2773
rect 218763 2745 218791 2773
rect 218577 876 218605 904
rect 218639 876 218667 904
rect 218701 876 218729 904
rect 218763 876 218791 904
rect 218577 814 218605 842
rect 218639 814 218667 842
rect 218701 814 218729 842
rect 218763 814 218791 842
rect 218577 752 218605 780
rect 218639 752 218667 780
rect 218701 752 218729 780
rect 218763 752 218791 780
rect 218577 690 218605 718
rect 218639 690 218667 718
rect 218701 690 218729 718
rect 218763 690 218791 718
rect 220437 5931 220465 5959
rect 220499 5931 220527 5959
rect 220561 5931 220589 5959
rect 220623 5931 220651 5959
rect 220437 5869 220465 5897
rect 220499 5869 220527 5897
rect 220561 5869 220589 5897
rect 220623 5869 220651 5897
rect 220437 5807 220465 5835
rect 220499 5807 220527 5835
rect 220561 5807 220589 5835
rect 220623 5807 220651 5835
rect 220437 5745 220465 5773
rect 220499 5745 220527 5773
rect 220561 5745 220589 5773
rect 220623 5745 220651 5773
rect 220437 396 220465 424
rect 220499 396 220527 424
rect 220561 396 220589 424
rect 220623 396 220651 424
rect 220437 334 220465 362
rect 220499 334 220527 362
rect 220561 334 220589 362
rect 220623 334 220651 362
rect 220437 272 220465 300
rect 220499 272 220527 300
rect 220561 272 220589 300
rect 220623 272 220651 300
rect 220437 210 220465 238
rect 220499 210 220527 238
rect 220561 210 220589 238
rect 220623 210 220651 238
rect 227577 11931 227605 11959
rect 227639 11931 227667 11959
rect 227701 11931 227729 11959
rect 227763 11931 227791 11959
rect 227577 11869 227605 11897
rect 227639 11869 227667 11897
rect 227701 11869 227729 11897
rect 227763 11869 227791 11897
rect 227577 11807 227605 11835
rect 227639 11807 227667 11835
rect 227701 11807 227729 11835
rect 227763 11807 227791 11835
rect 227577 11745 227605 11773
rect 227639 11745 227667 11773
rect 227701 11745 227729 11773
rect 227763 11745 227791 11773
rect 227577 2931 227605 2959
rect 227639 2931 227667 2959
rect 227701 2931 227729 2959
rect 227763 2931 227791 2959
rect 227577 2869 227605 2897
rect 227639 2869 227667 2897
rect 227701 2869 227729 2897
rect 227763 2869 227791 2897
rect 227577 2807 227605 2835
rect 227639 2807 227667 2835
rect 227701 2807 227729 2835
rect 227763 2807 227791 2835
rect 227577 2745 227605 2773
rect 227639 2745 227667 2773
rect 227701 2745 227729 2773
rect 227763 2745 227791 2773
rect 227577 876 227605 904
rect 227639 876 227667 904
rect 227701 876 227729 904
rect 227763 876 227791 904
rect 227577 814 227605 842
rect 227639 814 227667 842
rect 227701 814 227729 842
rect 227763 814 227791 842
rect 227577 752 227605 780
rect 227639 752 227667 780
rect 227701 752 227729 780
rect 227763 752 227791 780
rect 227577 690 227605 718
rect 227639 690 227667 718
rect 227701 690 227729 718
rect 227763 690 227791 718
rect 229437 5931 229465 5959
rect 229499 5931 229527 5959
rect 229561 5931 229589 5959
rect 229623 5931 229651 5959
rect 229437 5869 229465 5897
rect 229499 5869 229527 5897
rect 229561 5869 229589 5897
rect 229623 5869 229651 5897
rect 229437 5807 229465 5835
rect 229499 5807 229527 5835
rect 229561 5807 229589 5835
rect 229623 5807 229651 5835
rect 229437 5745 229465 5773
rect 229499 5745 229527 5773
rect 229561 5745 229589 5773
rect 229623 5745 229651 5773
rect 229437 396 229465 424
rect 229499 396 229527 424
rect 229561 396 229589 424
rect 229623 396 229651 424
rect 229437 334 229465 362
rect 229499 334 229527 362
rect 229561 334 229589 362
rect 229623 334 229651 362
rect 229437 272 229465 300
rect 229499 272 229527 300
rect 229561 272 229589 300
rect 229623 272 229651 300
rect 229437 210 229465 238
rect 229499 210 229527 238
rect 229561 210 229589 238
rect 229623 210 229651 238
rect 236577 11931 236605 11959
rect 236639 11931 236667 11959
rect 236701 11931 236729 11959
rect 236763 11931 236791 11959
rect 236577 11869 236605 11897
rect 236639 11869 236667 11897
rect 236701 11869 236729 11897
rect 236763 11869 236791 11897
rect 236577 11807 236605 11835
rect 236639 11807 236667 11835
rect 236701 11807 236729 11835
rect 236763 11807 236791 11835
rect 236577 11745 236605 11773
rect 236639 11745 236667 11773
rect 236701 11745 236729 11773
rect 236763 11745 236791 11773
rect 236577 2931 236605 2959
rect 236639 2931 236667 2959
rect 236701 2931 236729 2959
rect 236763 2931 236791 2959
rect 236577 2869 236605 2897
rect 236639 2869 236667 2897
rect 236701 2869 236729 2897
rect 236763 2869 236791 2897
rect 236577 2807 236605 2835
rect 236639 2807 236667 2835
rect 236701 2807 236729 2835
rect 236763 2807 236791 2835
rect 236577 2745 236605 2773
rect 236639 2745 236667 2773
rect 236701 2745 236729 2773
rect 236763 2745 236791 2773
rect 236577 876 236605 904
rect 236639 876 236667 904
rect 236701 876 236729 904
rect 236763 876 236791 904
rect 236577 814 236605 842
rect 236639 814 236667 842
rect 236701 814 236729 842
rect 236763 814 236791 842
rect 236577 752 236605 780
rect 236639 752 236667 780
rect 236701 752 236729 780
rect 236763 752 236791 780
rect 236577 690 236605 718
rect 236639 690 236667 718
rect 236701 690 236729 718
rect 236763 690 236791 718
rect 238437 5931 238465 5959
rect 238499 5931 238527 5959
rect 238561 5931 238589 5959
rect 238623 5931 238651 5959
rect 238437 5869 238465 5897
rect 238499 5869 238527 5897
rect 238561 5869 238589 5897
rect 238623 5869 238651 5897
rect 238437 5807 238465 5835
rect 238499 5807 238527 5835
rect 238561 5807 238589 5835
rect 238623 5807 238651 5835
rect 238437 5745 238465 5773
rect 238499 5745 238527 5773
rect 238561 5745 238589 5773
rect 238623 5745 238651 5773
rect 238437 396 238465 424
rect 238499 396 238527 424
rect 238561 396 238589 424
rect 238623 396 238651 424
rect 238437 334 238465 362
rect 238499 334 238527 362
rect 238561 334 238589 362
rect 238623 334 238651 362
rect 238437 272 238465 300
rect 238499 272 238527 300
rect 238561 272 238589 300
rect 238623 272 238651 300
rect 238437 210 238465 238
rect 238499 210 238527 238
rect 238561 210 238589 238
rect 238623 210 238651 238
rect 245577 11931 245605 11959
rect 245639 11931 245667 11959
rect 245701 11931 245729 11959
rect 245763 11931 245791 11959
rect 245577 11869 245605 11897
rect 245639 11869 245667 11897
rect 245701 11869 245729 11897
rect 245763 11869 245791 11897
rect 245577 11807 245605 11835
rect 245639 11807 245667 11835
rect 245701 11807 245729 11835
rect 245763 11807 245791 11835
rect 245577 11745 245605 11773
rect 245639 11745 245667 11773
rect 245701 11745 245729 11773
rect 245763 11745 245791 11773
rect 245577 2931 245605 2959
rect 245639 2931 245667 2959
rect 245701 2931 245729 2959
rect 245763 2931 245791 2959
rect 245577 2869 245605 2897
rect 245639 2869 245667 2897
rect 245701 2869 245729 2897
rect 245763 2869 245791 2897
rect 245577 2807 245605 2835
rect 245639 2807 245667 2835
rect 245701 2807 245729 2835
rect 245763 2807 245791 2835
rect 245577 2745 245605 2773
rect 245639 2745 245667 2773
rect 245701 2745 245729 2773
rect 245763 2745 245791 2773
rect 245577 876 245605 904
rect 245639 876 245667 904
rect 245701 876 245729 904
rect 245763 876 245791 904
rect 245577 814 245605 842
rect 245639 814 245667 842
rect 245701 814 245729 842
rect 245763 814 245791 842
rect 245577 752 245605 780
rect 245639 752 245667 780
rect 245701 752 245729 780
rect 245763 752 245791 780
rect 245577 690 245605 718
rect 245639 690 245667 718
rect 245701 690 245729 718
rect 245763 690 245791 718
rect 247437 5931 247465 5959
rect 247499 5931 247527 5959
rect 247561 5931 247589 5959
rect 247623 5931 247651 5959
rect 247437 5869 247465 5897
rect 247499 5869 247527 5897
rect 247561 5869 247589 5897
rect 247623 5869 247651 5897
rect 247437 5807 247465 5835
rect 247499 5807 247527 5835
rect 247561 5807 247589 5835
rect 247623 5807 247651 5835
rect 247437 5745 247465 5773
rect 247499 5745 247527 5773
rect 247561 5745 247589 5773
rect 247623 5745 247651 5773
rect 247437 396 247465 424
rect 247499 396 247527 424
rect 247561 396 247589 424
rect 247623 396 247651 424
rect 247437 334 247465 362
rect 247499 334 247527 362
rect 247561 334 247589 362
rect 247623 334 247651 362
rect 247437 272 247465 300
rect 247499 272 247527 300
rect 247561 272 247589 300
rect 247623 272 247651 300
rect 247437 210 247465 238
rect 247499 210 247527 238
rect 247561 210 247589 238
rect 247623 210 247651 238
rect 256437 248931 256465 248959
rect 256499 248931 256527 248959
rect 256561 248931 256589 248959
rect 256623 248931 256651 248959
rect 256437 248869 256465 248897
rect 256499 248869 256527 248897
rect 256561 248869 256589 248897
rect 256623 248869 256651 248897
rect 256437 248807 256465 248835
rect 256499 248807 256527 248835
rect 256561 248807 256589 248835
rect 256623 248807 256651 248835
rect 256437 248745 256465 248773
rect 256499 248745 256527 248773
rect 256561 248745 256589 248773
rect 256623 248745 256651 248773
rect 256437 239931 256465 239959
rect 256499 239931 256527 239959
rect 256561 239931 256589 239959
rect 256623 239931 256651 239959
rect 256437 239869 256465 239897
rect 256499 239869 256527 239897
rect 256561 239869 256589 239897
rect 256623 239869 256651 239897
rect 256437 239807 256465 239835
rect 256499 239807 256527 239835
rect 256561 239807 256589 239835
rect 256623 239807 256651 239835
rect 256437 239745 256465 239773
rect 256499 239745 256527 239773
rect 256561 239745 256589 239773
rect 256623 239745 256651 239773
rect 256437 230931 256465 230959
rect 256499 230931 256527 230959
rect 256561 230931 256589 230959
rect 256623 230931 256651 230959
rect 256437 230869 256465 230897
rect 256499 230869 256527 230897
rect 256561 230869 256589 230897
rect 256623 230869 256651 230897
rect 256437 230807 256465 230835
rect 256499 230807 256527 230835
rect 256561 230807 256589 230835
rect 256623 230807 256651 230835
rect 256437 230745 256465 230773
rect 256499 230745 256527 230773
rect 256561 230745 256589 230773
rect 256623 230745 256651 230773
rect 256437 221931 256465 221959
rect 256499 221931 256527 221959
rect 256561 221931 256589 221959
rect 256623 221931 256651 221959
rect 256437 221869 256465 221897
rect 256499 221869 256527 221897
rect 256561 221869 256589 221897
rect 256623 221869 256651 221897
rect 256437 221807 256465 221835
rect 256499 221807 256527 221835
rect 256561 221807 256589 221835
rect 256623 221807 256651 221835
rect 256437 221745 256465 221773
rect 256499 221745 256527 221773
rect 256561 221745 256589 221773
rect 256623 221745 256651 221773
rect 256437 212931 256465 212959
rect 256499 212931 256527 212959
rect 256561 212931 256589 212959
rect 256623 212931 256651 212959
rect 256437 212869 256465 212897
rect 256499 212869 256527 212897
rect 256561 212869 256589 212897
rect 256623 212869 256651 212897
rect 256437 212807 256465 212835
rect 256499 212807 256527 212835
rect 256561 212807 256589 212835
rect 256623 212807 256651 212835
rect 256437 212745 256465 212773
rect 256499 212745 256527 212773
rect 256561 212745 256589 212773
rect 256623 212745 256651 212773
rect 256437 203931 256465 203959
rect 256499 203931 256527 203959
rect 256561 203931 256589 203959
rect 256623 203931 256651 203959
rect 256437 203869 256465 203897
rect 256499 203869 256527 203897
rect 256561 203869 256589 203897
rect 256623 203869 256651 203897
rect 256437 203807 256465 203835
rect 256499 203807 256527 203835
rect 256561 203807 256589 203835
rect 256623 203807 256651 203835
rect 256437 203745 256465 203773
rect 256499 203745 256527 203773
rect 256561 203745 256589 203773
rect 256623 203745 256651 203773
rect 256437 194931 256465 194959
rect 256499 194931 256527 194959
rect 256561 194931 256589 194959
rect 256623 194931 256651 194959
rect 256437 194869 256465 194897
rect 256499 194869 256527 194897
rect 256561 194869 256589 194897
rect 256623 194869 256651 194897
rect 256437 194807 256465 194835
rect 256499 194807 256527 194835
rect 256561 194807 256589 194835
rect 256623 194807 256651 194835
rect 256437 194745 256465 194773
rect 256499 194745 256527 194773
rect 256561 194745 256589 194773
rect 256623 194745 256651 194773
rect 256437 185931 256465 185959
rect 256499 185931 256527 185959
rect 256561 185931 256589 185959
rect 256623 185931 256651 185959
rect 256437 185869 256465 185897
rect 256499 185869 256527 185897
rect 256561 185869 256589 185897
rect 256623 185869 256651 185897
rect 256437 185807 256465 185835
rect 256499 185807 256527 185835
rect 256561 185807 256589 185835
rect 256623 185807 256651 185835
rect 256437 185745 256465 185773
rect 256499 185745 256527 185773
rect 256561 185745 256589 185773
rect 256623 185745 256651 185773
rect 256437 176931 256465 176959
rect 256499 176931 256527 176959
rect 256561 176931 256589 176959
rect 256623 176931 256651 176959
rect 256437 176869 256465 176897
rect 256499 176869 256527 176897
rect 256561 176869 256589 176897
rect 256623 176869 256651 176897
rect 256437 176807 256465 176835
rect 256499 176807 256527 176835
rect 256561 176807 256589 176835
rect 256623 176807 256651 176835
rect 256437 176745 256465 176773
rect 256499 176745 256527 176773
rect 256561 176745 256589 176773
rect 256623 176745 256651 176773
rect 256437 167931 256465 167959
rect 256499 167931 256527 167959
rect 256561 167931 256589 167959
rect 256623 167931 256651 167959
rect 256437 167869 256465 167897
rect 256499 167869 256527 167897
rect 256561 167869 256589 167897
rect 256623 167869 256651 167897
rect 256437 167807 256465 167835
rect 256499 167807 256527 167835
rect 256561 167807 256589 167835
rect 256623 167807 256651 167835
rect 256437 167745 256465 167773
rect 256499 167745 256527 167773
rect 256561 167745 256589 167773
rect 256623 167745 256651 167773
rect 256437 158931 256465 158959
rect 256499 158931 256527 158959
rect 256561 158931 256589 158959
rect 256623 158931 256651 158959
rect 256437 158869 256465 158897
rect 256499 158869 256527 158897
rect 256561 158869 256589 158897
rect 256623 158869 256651 158897
rect 256437 158807 256465 158835
rect 256499 158807 256527 158835
rect 256561 158807 256589 158835
rect 256623 158807 256651 158835
rect 256437 158745 256465 158773
rect 256499 158745 256527 158773
rect 256561 158745 256589 158773
rect 256623 158745 256651 158773
rect 256437 149931 256465 149959
rect 256499 149931 256527 149959
rect 256561 149931 256589 149959
rect 256623 149931 256651 149959
rect 256437 149869 256465 149897
rect 256499 149869 256527 149897
rect 256561 149869 256589 149897
rect 256623 149869 256651 149897
rect 256437 149807 256465 149835
rect 256499 149807 256527 149835
rect 256561 149807 256589 149835
rect 256623 149807 256651 149835
rect 256437 149745 256465 149773
rect 256499 149745 256527 149773
rect 256561 149745 256589 149773
rect 256623 149745 256651 149773
rect 256437 140931 256465 140959
rect 256499 140931 256527 140959
rect 256561 140931 256589 140959
rect 256623 140931 256651 140959
rect 256437 140869 256465 140897
rect 256499 140869 256527 140897
rect 256561 140869 256589 140897
rect 256623 140869 256651 140897
rect 256437 140807 256465 140835
rect 256499 140807 256527 140835
rect 256561 140807 256589 140835
rect 256623 140807 256651 140835
rect 256437 140745 256465 140773
rect 256499 140745 256527 140773
rect 256561 140745 256589 140773
rect 256623 140745 256651 140773
rect 256437 131931 256465 131959
rect 256499 131931 256527 131959
rect 256561 131931 256589 131959
rect 256623 131931 256651 131959
rect 256437 131869 256465 131897
rect 256499 131869 256527 131897
rect 256561 131869 256589 131897
rect 256623 131869 256651 131897
rect 256437 131807 256465 131835
rect 256499 131807 256527 131835
rect 256561 131807 256589 131835
rect 256623 131807 256651 131835
rect 256437 131745 256465 131773
rect 256499 131745 256527 131773
rect 256561 131745 256589 131773
rect 256623 131745 256651 131773
rect 256437 122931 256465 122959
rect 256499 122931 256527 122959
rect 256561 122931 256589 122959
rect 256623 122931 256651 122959
rect 256437 122869 256465 122897
rect 256499 122869 256527 122897
rect 256561 122869 256589 122897
rect 256623 122869 256651 122897
rect 256437 122807 256465 122835
rect 256499 122807 256527 122835
rect 256561 122807 256589 122835
rect 256623 122807 256651 122835
rect 256437 122745 256465 122773
rect 256499 122745 256527 122773
rect 256561 122745 256589 122773
rect 256623 122745 256651 122773
rect 256437 113931 256465 113959
rect 256499 113931 256527 113959
rect 256561 113931 256589 113959
rect 256623 113931 256651 113959
rect 256437 113869 256465 113897
rect 256499 113869 256527 113897
rect 256561 113869 256589 113897
rect 256623 113869 256651 113897
rect 256437 113807 256465 113835
rect 256499 113807 256527 113835
rect 256561 113807 256589 113835
rect 256623 113807 256651 113835
rect 256437 113745 256465 113773
rect 256499 113745 256527 113773
rect 256561 113745 256589 113773
rect 256623 113745 256651 113773
rect 256437 104931 256465 104959
rect 256499 104931 256527 104959
rect 256561 104931 256589 104959
rect 256623 104931 256651 104959
rect 256437 104869 256465 104897
rect 256499 104869 256527 104897
rect 256561 104869 256589 104897
rect 256623 104869 256651 104897
rect 256437 104807 256465 104835
rect 256499 104807 256527 104835
rect 256561 104807 256589 104835
rect 256623 104807 256651 104835
rect 256437 104745 256465 104773
rect 256499 104745 256527 104773
rect 256561 104745 256589 104773
rect 256623 104745 256651 104773
rect 256437 95931 256465 95959
rect 256499 95931 256527 95959
rect 256561 95931 256589 95959
rect 256623 95931 256651 95959
rect 256437 95869 256465 95897
rect 256499 95869 256527 95897
rect 256561 95869 256589 95897
rect 256623 95869 256651 95897
rect 256437 95807 256465 95835
rect 256499 95807 256527 95835
rect 256561 95807 256589 95835
rect 256623 95807 256651 95835
rect 256437 95745 256465 95773
rect 256499 95745 256527 95773
rect 256561 95745 256589 95773
rect 256623 95745 256651 95773
rect 256437 86931 256465 86959
rect 256499 86931 256527 86959
rect 256561 86931 256589 86959
rect 256623 86931 256651 86959
rect 256437 86869 256465 86897
rect 256499 86869 256527 86897
rect 256561 86869 256589 86897
rect 256623 86869 256651 86897
rect 256437 86807 256465 86835
rect 256499 86807 256527 86835
rect 256561 86807 256589 86835
rect 256623 86807 256651 86835
rect 256437 86745 256465 86773
rect 256499 86745 256527 86773
rect 256561 86745 256589 86773
rect 256623 86745 256651 86773
rect 256437 77931 256465 77959
rect 256499 77931 256527 77959
rect 256561 77931 256589 77959
rect 256623 77931 256651 77959
rect 256437 77869 256465 77897
rect 256499 77869 256527 77897
rect 256561 77869 256589 77897
rect 256623 77869 256651 77897
rect 256437 77807 256465 77835
rect 256499 77807 256527 77835
rect 256561 77807 256589 77835
rect 256623 77807 256651 77835
rect 256437 77745 256465 77773
rect 256499 77745 256527 77773
rect 256561 77745 256589 77773
rect 256623 77745 256651 77773
rect 256437 68931 256465 68959
rect 256499 68931 256527 68959
rect 256561 68931 256589 68959
rect 256623 68931 256651 68959
rect 256437 68869 256465 68897
rect 256499 68869 256527 68897
rect 256561 68869 256589 68897
rect 256623 68869 256651 68897
rect 256437 68807 256465 68835
rect 256499 68807 256527 68835
rect 256561 68807 256589 68835
rect 256623 68807 256651 68835
rect 256437 68745 256465 68773
rect 256499 68745 256527 68773
rect 256561 68745 256589 68773
rect 256623 68745 256651 68773
rect 256437 59931 256465 59959
rect 256499 59931 256527 59959
rect 256561 59931 256589 59959
rect 256623 59931 256651 59959
rect 256437 59869 256465 59897
rect 256499 59869 256527 59897
rect 256561 59869 256589 59897
rect 256623 59869 256651 59897
rect 256437 59807 256465 59835
rect 256499 59807 256527 59835
rect 256561 59807 256589 59835
rect 256623 59807 256651 59835
rect 256437 59745 256465 59773
rect 256499 59745 256527 59773
rect 256561 59745 256589 59773
rect 256623 59745 256651 59773
rect 256437 50931 256465 50959
rect 256499 50931 256527 50959
rect 256561 50931 256589 50959
rect 256623 50931 256651 50959
rect 256437 50869 256465 50897
rect 256499 50869 256527 50897
rect 256561 50869 256589 50897
rect 256623 50869 256651 50897
rect 256437 50807 256465 50835
rect 256499 50807 256527 50835
rect 256561 50807 256589 50835
rect 256623 50807 256651 50835
rect 256437 50745 256465 50773
rect 256499 50745 256527 50773
rect 256561 50745 256589 50773
rect 256623 50745 256651 50773
rect 256437 41931 256465 41959
rect 256499 41931 256527 41959
rect 256561 41931 256589 41959
rect 256623 41931 256651 41959
rect 256437 41869 256465 41897
rect 256499 41869 256527 41897
rect 256561 41869 256589 41897
rect 256623 41869 256651 41897
rect 256437 41807 256465 41835
rect 256499 41807 256527 41835
rect 256561 41807 256589 41835
rect 256623 41807 256651 41835
rect 256437 41745 256465 41773
rect 256499 41745 256527 41773
rect 256561 41745 256589 41773
rect 256623 41745 256651 41773
rect 256437 32931 256465 32959
rect 256499 32931 256527 32959
rect 256561 32931 256589 32959
rect 256623 32931 256651 32959
rect 256437 32869 256465 32897
rect 256499 32869 256527 32897
rect 256561 32869 256589 32897
rect 256623 32869 256651 32897
rect 256437 32807 256465 32835
rect 256499 32807 256527 32835
rect 256561 32807 256589 32835
rect 256623 32807 256651 32835
rect 256437 32745 256465 32773
rect 256499 32745 256527 32773
rect 256561 32745 256589 32773
rect 256623 32745 256651 32773
rect 256437 23931 256465 23959
rect 256499 23931 256527 23959
rect 256561 23931 256589 23959
rect 256623 23931 256651 23959
rect 256437 23869 256465 23897
rect 256499 23869 256527 23897
rect 256561 23869 256589 23897
rect 256623 23869 256651 23897
rect 256437 23807 256465 23835
rect 256499 23807 256527 23835
rect 256561 23807 256589 23835
rect 256623 23807 256651 23835
rect 256437 23745 256465 23773
rect 256499 23745 256527 23773
rect 256561 23745 256589 23773
rect 256623 23745 256651 23773
rect 256437 14931 256465 14959
rect 256499 14931 256527 14959
rect 256561 14931 256589 14959
rect 256623 14931 256651 14959
rect 256437 14869 256465 14897
rect 256499 14869 256527 14897
rect 256561 14869 256589 14897
rect 256623 14869 256651 14897
rect 256437 14807 256465 14835
rect 256499 14807 256527 14835
rect 256561 14807 256589 14835
rect 256623 14807 256651 14835
rect 256437 14745 256465 14773
rect 256499 14745 256527 14773
rect 256561 14745 256589 14773
rect 256623 14745 256651 14773
rect 254577 11931 254605 11959
rect 254639 11931 254667 11959
rect 254701 11931 254729 11959
rect 254763 11931 254791 11959
rect 254577 11869 254605 11897
rect 254639 11869 254667 11897
rect 254701 11869 254729 11897
rect 254763 11869 254791 11897
rect 254577 11807 254605 11835
rect 254639 11807 254667 11835
rect 254701 11807 254729 11835
rect 254763 11807 254791 11835
rect 254577 11745 254605 11773
rect 254639 11745 254667 11773
rect 254701 11745 254729 11773
rect 254763 11745 254791 11773
rect 254577 2931 254605 2959
rect 254639 2931 254667 2959
rect 254701 2931 254729 2959
rect 254763 2931 254791 2959
rect 254577 2869 254605 2897
rect 254639 2869 254667 2897
rect 254701 2869 254729 2897
rect 254763 2869 254791 2897
rect 254577 2807 254605 2835
rect 254639 2807 254667 2835
rect 254701 2807 254729 2835
rect 254763 2807 254791 2835
rect 254577 2745 254605 2773
rect 254639 2745 254667 2773
rect 254701 2745 254729 2773
rect 254763 2745 254791 2773
rect 254577 876 254605 904
rect 254639 876 254667 904
rect 254701 876 254729 904
rect 254763 876 254791 904
rect 254577 814 254605 842
rect 254639 814 254667 842
rect 254701 814 254729 842
rect 254763 814 254791 842
rect 254577 752 254605 780
rect 254639 752 254667 780
rect 254701 752 254729 780
rect 254763 752 254791 780
rect 254577 690 254605 718
rect 254639 690 254667 718
rect 254701 690 254729 718
rect 254763 690 254791 718
rect 256437 5931 256465 5959
rect 256499 5931 256527 5959
rect 256561 5931 256589 5959
rect 256623 5931 256651 5959
rect 256437 5869 256465 5897
rect 256499 5869 256527 5897
rect 256561 5869 256589 5897
rect 256623 5869 256651 5897
rect 256437 5807 256465 5835
rect 256499 5807 256527 5835
rect 256561 5807 256589 5835
rect 256623 5807 256651 5835
rect 256437 5745 256465 5773
rect 256499 5745 256527 5773
rect 256561 5745 256589 5773
rect 256623 5745 256651 5773
rect 256437 396 256465 424
rect 256499 396 256527 424
rect 256561 396 256589 424
rect 256623 396 256651 424
rect 256437 334 256465 362
rect 256499 334 256527 362
rect 256561 334 256589 362
rect 256623 334 256651 362
rect 256437 272 256465 300
rect 256499 272 256527 300
rect 256561 272 256589 300
rect 256623 272 256651 300
rect 256437 210 256465 238
rect 256499 210 256527 238
rect 256561 210 256589 238
rect 256623 210 256651 238
rect 263577 299162 263605 299190
rect 263639 299162 263667 299190
rect 263701 299162 263729 299190
rect 263763 299162 263791 299190
rect 263577 299100 263605 299128
rect 263639 299100 263667 299128
rect 263701 299100 263729 299128
rect 263763 299100 263791 299128
rect 263577 299038 263605 299066
rect 263639 299038 263667 299066
rect 263701 299038 263729 299066
rect 263763 299038 263791 299066
rect 263577 298976 263605 299004
rect 263639 298976 263667 299004
rect 263701 298976 263729 299004
rect 263763 298976 263791 299004
rect 263577 290931 263605 290959
rect 263639 290931 263667 290959
rect 263701 290931 263729 290959
rect 263763 290931 263791 290959
rect 263577 290869 263605 290897
rect 263639 290869 263667 290897
rect 263701 290869 263729 290897
rect 263763 290869 263791 290897
rect 263577 290807 263605 290835
rect 263639 290807 263667 290835
rect 263701 290807 263729 290835
rect 263763 290807 263791 290835
rect 263577 290745 263605 290773
rect 263639 290745 263667 290773
rect 263701 290745 263729 290773
rect 263763 290745 263791 290773
rect 263577 281931 263605 281959
rect 263639 281931 263667 281959
rect 263701 281931 263729 281959
rect 263763 281931 263791 281959
rect 263577 281869 263605 281897
rect 263639 281869 263667 281897
rect 263701 281869 263729 281897
rect 263763 281869 263791 281897
rect 263577 281807 263605 281835
rect 263639 281807 263667 281835
rect 263701 281807 263729 281835
rect 263763 281807 263791 281835
rect 263577 281745 263605 281773
rect 263639 281745 263667 281773
rect 263701 281745 263729 281773
rect 263763 281745 263791 281773
rect 263577 272931 263605 272959
rect 263639 272931 263667 272959
rect 263701 272931 263729 272959
rect 263763 272931 263791 272959
rect 263577 272869 263605 272897
rect 263639 272869 263667 272897
rect 263701 272869 263729 272897
rect 263763 272869 263791 272897
rect 263577 272807 263605 272835
rect 263639 272807 263667 272835
rect 263701 272807 263729 272835
rect 263763 272807 263791 272835
rect 263577 272745 263605 272773
rect 263639 272745 263667 272773
rect 263701 272745 263729 272773
rect 263763 272745 263791 272773
rect 263577 263931 263605 263959
rect 263639 263931 263667 263959
rect 263701 263931 263729 263959
rect 263763 263931 263791 263959
rect 263577 263869 263605 263897
rect 263639 263869 263667 263897
rect 263701 263869 263729 263897
rect 263763 263869 263791 263897
rect 263577 263807 263605 263835
rect 263639 263807 263667 263835
rect 263701 263807 263729 263835
rect 263763 263807 263791 263835
rect 263577 263745 263605 263773
rect 263639 263745 263667 263773
rect 263701 263745 263729 263773
rect 263763 263745 263791 263773
rect 263577 254931 263605 254959
rect 263639 254931 263667 254959
rect 263701 254931 263729 254959
rect 263763 254931 263791 254959
rect 263577 254869 263605 254897
rect 263639 254869 263667 254897
rect 263701 254869 263729 254897
rect 263763 254869 263791 254897
rect 263577 254807 263605 254835
rect 263639 254807 263667 254835
rect 263701 254807 263729 254835
rect 263763 254807 263791 254835
rect 263577 254745 263605 254773
rect 263639 254745 263667 254773
rect 263701 254745 263729 254773
rect 263763 254745 263791 254773
rect 263577 245931 263605 245959
rect 263639 245931 263667 245959
rect 263701 245931 263729 245959
rect 263763 245931 263791 245959
rect 263577 245869 263605 245897
rect 263639 245869 263667 245897
rect 263701 245869 263729 245897
rect 263763 245869 263791 245897
rect 263577 245807 263605 245835
rect 263639 245807 263667 245835
rect 263701 245807 263729 245835
rect 263763 245807 263791 245835
rect 263577 245745 263605 245773
rect 263639 245745 263667 245773
rect 263701 245745 263729 245773
rect 263763 245745 263791 245773
rect 263577 236931 263605 236959
rect 263639 236931 263667 236959
rect 263701 236931 263729 236959
rect 263763 236931 263791 236959
rect 263577 236869 263605 236897
rect 263639 236869 263667 236897
rect 263701 236869 263729 236897
rect 263763 236869 263791 236897
rect 263577 236807 263605 236835
rect 263639 236807 263667 236835
rect 263701 236807 263729 236835
rect 263763 236807 263791 236835
rect 263577 236745 263605 236773
rect 263639 236745 263667 236773
rect 263701 236745 263729 236773
rect 263763 236745 263791 236773
rect 263577 227931 263605 227959
rect 263639 227931 263667 227959
rect 263701 227931 263729 227959
rect 263763 227931 263791 227959
rect 263577 227869 263605 227897
rect 263639 227869 263667 227897
rect 263701 227869 263729 227897
rect 263763 227869 263791 227897
rect 263577 227807 263605 227835
rect 263639 227807 263667 227835
rect 263701 227807 263729 227835
rect 263763 227807 263791 227835
rect 263577 227745 263605 227773
rect 263639 227745 263667 227773
rect 263701 227745 263729 227773
rect 263763 227745 263791 227773
rect 263577 218931 263605 218959
rect 263639 218931 263667 218959
rect 263701 218931 263729 218959
rect 263763 218931 263791 218959
rect 263577 218869 263605 218897
rect 263639 218869 263667 218897
rect 263701 218869 263729 218897
rect 263763 218869 263791 218897
rect 263577 218807 263605 218835
rect 263639 218807 263667 218835
rect 263701 218807 263729 218835
rect 263763 218807 263791 218835
rect 263577 218745 263605 218773
rect 263639 218745 263667 218773
rect 263701 218745 263729 218773
rect 263763 218745 263791 218773
rect 263577 209931 263605 209959
rect 263639 209931 263667 209959
rect 263701 209931 263729 209959
rect 263763 209931 263791 209959
rect 263577 209869 263605 209897
rect 263639 209869 263667 209897
rect 263701 209869 263729 209897
rect 263763 209869 263791 209897
rect 263577 209807 263605 209835
rect 263639 209807 263667 209835
rect 263701 209807 263729 209835
rect 263763 209807 263791 209835
rect 263577 209745 263605 209773
rect 263639 209745 263667 209773
rect 263701 209745 263729 209773
rect 263763 209745 263791 209773
rect 263577 200931 263605 200959
rect 263639 200931 263667 200959
rect 263701 200931 263729 200959
rect 263763 200931 263791 200959
rect 263577 200869 263605 200897
rect 263639 200869 263667 200897
rect 263701 200869 263729 200897
rect 263763 200869 263791 200897
rect 263577 200807 263605 200835
rect 263639 200807 263667 200835
rect 263701 200807 263729 200835
rect 263763 200807 263791 200835
rect 263577 200745 263605 200773
rect 263639 200745 263667 200773
rect 263701 200745 263729 200773
rect 263763 200745 263791 200773
rect 263577 191931 263605 191959
rect 263639 191931 263667 191959
rect 263701 191931 263729 191959
rect 263763 191931 263791 191959
rect 263577 191869 263605 191897
rect 263639 191869 263667 191897
rect 263701 191869 263729 191897
rect 263763 191869 263791 191897
rect 263577 191807 263605 191835
rect 263639 191807 263667 191835
rect 263701 191807 263729 191835
rect 263763 191807 263791 191835
rect 263577 191745 263605 191773
rect 263639 191745 263667 191773
rect 263701 191745 263729 191773
rect 263763 191745 263791 191773
rect 263577 182931 263605 182959
rect 263639 182931 263667 182959
rect 263701 182931 263729 182959
rect 263763 182931 263791 182959
rect 263577 182869 263605 182897
rect 263639 182869 263667 182897
rect 263701 182869 263729 182897
rect 263763 182869 263791 182897
rect 263577 182807 263605 182835
rect 263639 182807 263667 182835
rect 263701 182807 263729 182835
rect 263763 182807 263791 182835
rect 263577 182745 263605 182773
rect 263639 182745 263667 182773
rect 263701 182745 263729 182773
rect 263763 182745 263791 182773
rect 263577 173931 263605 173959
rect 263639 173931 263667 173959
rect 263701 173931 263729 173959
rect 263763 173931 263791 173959
rect 263577 173869 263605 173897
rect 263639 173869 263667 173897
rect 263701 173869 263729 173897
rect 263763 173869 263791 173897
rect 263577 173807 263605 173835
rect 263639 173807 263667 173835
rect 263701 173807 263729 173835
rect 263763 173807 263791 173835
rect 263577 173745 263605 173773
rect 263639 173745 263667 173773
rect 263701 173745 263729 173773
rect 263763 173745 263791 173773
rect 263577 164931 263605 164959
rect 263639 164931 263667 164959
rect 263701 164931 263729 164959
rect 263763 164931 263791 164959
rect 263577 164869 263605 164897
rect 263639 164869 263667 164897
rect 263701 164869 263729 164897
rect 263763 164869 263791 164897
rect 263577 164807 263605 164835
rect 263639 164807 263667 164835
rect 263701 164807 263729 164835
rect 263763 164807 263791 164835
rect 263577 164745 263605 164773
rect 263639 164745 263667 164773
rect 263701 164745 263729 164773
rect 263763 164745 263791 164773
rect 263577 155931 263605 155959
rect 263639 155931 263667 155959
rect 263701 155931 263729 155959
rect 263763 155931 263791 155959
rect 263577 155869 263605 155897
rect 263639 155869 263667 155897
rect 263701 155869 263729 155897
rect 263763 155869 263791 155897
rect 263577 155807 263605 155835
rect 263639 155807 263667 155835
rect 263701 155807 263729 155835
rect 263763 155807 263791 155835
rect 263577 155745 263605 155773
rect 263639 155745 263667 155773
rect 263701 155745 263729 155773
rect 263763 155745 263791 155773
rect 263577 146931 263605 146959
rect 263639 146931 263667 146959
rect 263701 146931 263729 146959
rect 263763 146931 263791 146959
rect 263577 146869 263605 146897
rect 263639 146869 263667 146897
rect 263701 146869 263729 146897
rect 263763 146869 263791 146897
rect 263577 146807 263605 146835
rect 263639 146807 263667 146835
rect 263701 146807 263729 146835
rect 263763 146807 263791 146835
rect 263577 146745 263605 146773
rect 263639 146745 263667 146773
rect 263701 146745 263729 146773
rect 263763 146745 263791 146773
rect 263577 137931 263605 137959
rect 263639 137931 263667 137959
rect 263701 137931 263729 137959
rect 263763 137931 263791 137959
rect 263577 137869 263605 137897
rect 263639 137869 263667 137897
rect 263701 137869 263729 137897
rect 263763 137869 263791 137897
rect 263577 137807 263605 137835
rect 263639 137807 263667 137835
rect 263701 137807 263729 137835
rect 263763 137807 263791 137835
rect 263577 137745 263605 137773
rect 263639 137745 263667 137773
rect 263701 137745 263729 137773
rect 263763 137745 263791 137773
rect 263577 128931 263605 128959
rect 263639 128931 263667 128959
rect 263701 128931 263729 128959
rect 263763 128931 263791 128959
rect 263577 128869 263605 128897
rect 263639 128869 263667 128897
rect 263701 128869 263729 128897
rect 263763 128869 263791 128897
rect 263577 128807 263605 128835
rect 263639 128807 263667 128835
rect 263701 128807 263729 128835
rect 263763 128807 263791 128835
rect 263577 128745 263605 128773
rect 263639 128745 263667 128773
rect 263701 128745 263729 128773
rect 263763 128745 263791 128773
rect 263577 119931 263605 119959
rect 263639 119931 263667 119959
rect 263701 119931 263729 119959
rect 263763 119931 263791 119959
rect 263577 119869 263605 119897
rect 263639 119869 263667 119897
rect 263701 119869 263729 119897
rect 263763 119869 263791 119897
rect 263577 119807 263605 119835
rect 263639 119807 263667 119835
rect 263701 119807 263729 119835
rect 263763 119807 263791 119835
rect 263577 119745 263605 119773
rect 263639 119745 263667 119773
rect 263701 119745 263729 119773
rect 263763 119745 263791 119773
rect 263577 110931 263605 110959
rect 263639 110931 263667 110959
rect 263701 110931 263729 110959
rect 263763 110931 263791 110959
rect 263577 110869 263605 110897
rect 263639 110869 263667 110897
rect 263701 110869 263729 110897
rect 263763 110869 263791 110897
rect 263577 110807 263605 110835
rect 263639 110807 263667 110835
rect 263701 110807 263729 110835
rect 263763 110807 263791 110835
rect 263577 110745 263605 110773
rect 263639 110745 263667 110773
rect 263701 110745 263729 110773
rect 263763 110745 263791 110773
rect 263577 101931 263605 101959
rect 263639 101931 263667 101959
rect 263701 101931 263729 101959
rect 263763 101931 263791 101959
rect 263577 101869 263605 101897
rect 263639 101869 263667 101897
rect 263701 101869 263729 101897
rect 263763 101869 263791 101897
rect 263577 101807 263605 101835
rect 263639 101807 263667 101835
rect 263701 101807 263729 101835
rect 263763 101807 263791 101835
rect 263577 101745 263605 101773
rect 263639 101745 263667 101773
rect 263701 101745 263729 101773
rect 263763 101745 263791 101773
rect 263577 92931 263605 92959
rect 263639 92931 263667 92959
rect 263701 92931 263729 92959
rect 263763 92931 263791 92959
rect 263577 92869 263605 92897
rect 263639 92869 263667 92897
rect 263701 92869 263729 92897
rect 263763 92869 263791 92897
rect 263577 92807 263605 92835
rect 263639 92807 263667 92835
rect 263701 92807 263729 92835
rect 263763 92807 263791 92835
rect 263577 92745 263605 92773
rect 263639 92745 263667 92773
rect 263701 92745 263729 92773
rect 263763 92745 263791 92773
rect 263577 83931 263605 83959
rect 263639 83931 263667 83959
rect 263701 83931 263729 83959
rect 263763 83931 263791 83959
rect 263577 83869 263605 83897
rect 263639 83869 263667 83897
rect 263701 83869 263729 83897
rect 263763 83869 263791 83897
rect 263577 83807 263605 83835
rect 263639 83807 263667 83835
rect 263701 83807 263729 83835
rect 263763 83807 263791 83835
rect 263577 83745 263605 83773
rect 263639 83745 263667 83773
rect 263701 83745 263729 83773
rect 263763 83745 263791 83773
rect 263577 74931 263605 74959
rect 263639 74931 263667 74959
rect 263701 74931 263729 74959
rect 263763 74931 263791 74959
rect 263577 74869 263605 74897
rect 263639 74869 263667 74897
rect 263701 74869 263729 74897
rect 263763 74869 263791 74897
rect 263577 74807 263605 74835
rect 263639 74807 263667 74835
rect 263701 74807 263729 74835
rect 263763 74807 263791 74835
rect 263577 74745 263605 74773
rect 263639 74745 263667 74773
rect 263701 74745 263729 74773
rect 263763 74745 263791 74773
rect 263577 65931 263605 65959
rect 263639 65931 263667 65959
rect 263701 65931 263729 65959
rect 263763 65931 263791 65959
rect 263577 65869 263605 65897
rect 263639 65869 263667 65897
rect 263701 65869 263729 65897
rect 263763 65869 263791 65897
rect 263577 65807 263605 65835
rect 263639 65807 263667 65835
rect 263701 65807 263729 65835
rect 263763 65807 263791 65835
rect 263577 65745 263605 65773
rect 263639 65745 263667 65773
rect 263701 65745 263729 65773
rect 263763 65745 263791 65773
rect 263577 56931 263605 56959
rect 263639 56931 263667 56959
rect 263701 56931 263729 56959
rect 263763 56931 263791 56959
rect 263577 56869 263605 56897
rect 263639 56869 263667 56897
rect 263701 56869 263729 56897
rect 263763 56869 263791 56897
rect 263577 56807 263605 56835
rect 263639 56807 263667 56835
rect 263701 56807 263729 56835
rect 263763 56807 263791 56835
rect 263577 56745 263605 56773
rect 263639 56745 263667 56773
rect 263701 56745 263729 56773
rect 263763 56745 263791 56773
rect 263577 47931 263605 47959
rect 263639 47931 263667 47959
rect 263701 47931 263729 47959
rect 263763 47931 263791 47959
rect 263577 47869 263605 47897
rect 263639 47869 263667 47897
rect 263701 47869 263729 47897
rect 263763 47869 263791 47897
rect 263577 47807 263605 47835
rect 263639 47807 263667 47835
rect 263701 47807 263729 47835
rect 263763 47807 263791 47835
rect 263577 47745 263605 47773
rect 263639 47745 263667 47773
rect 263701 47745 263729 47773
rect 263763 47745 263791 47773
rect 263577 38931 263605 38959
rect 263639 38931 263667 38959
rect 263701 38931 263729 38959
rect 263763 38931 263791 38959
rect 263577 38869 263605 38897
rect 263639 38869 263667 38897
rect 263701 38869 263729 38897
rect 263763 38869 263791 38897
rect 263577 38807 263605 38835
rect 263639 38807 263667 38835
rect 263701 38807 263729 38835
rect 263763 38807 263791 38835
rect 263577 38745 263605 38773
rect 263639 38745 263667 38773
rect 263701 38745 263729 38773
rect 263763 38745 263791 38773
rect 263577 29931 263605 29959
rect 263639 29931 263667 29959
rect 263701 29931 263729 29959
rect 263763 29931 263791 29959
rect 263577 29869 263605 29897
rect 263639 29869 263667 29897
rect 263701 29869 263729 29897
rect 263763 29869 263791 29897
rect 263577 29807 263605 29835
rect 263639 29807 263667 29835
rect 263701 29807 263729 29835
rect 263763 29807 263791 29835
rect 263577 29745 263605 29773
rect 263639 29745 263667 29773
rect 263701 29745 263729 29773
rect 263763 29745 263791 29773
rect 263577 20931 263605 20959
rect 263639 20931 263667 20959
rect 263701 20931 263729 20959
rect 263763 20931 263791 20959
rect 263577 20869 263605 20897
rect 263639 20869 263667 20897
rect 263701 20869 263729 20897
rect 263763 20869 263791 20897
rect 263577 20807 263605 20835
rect 263639 20807 263667 20835
rect 263701 20807 263729 20835
rect 263763 20807 263791 20835
rect 263577 20745 263605 20773
rect 263639 20745 263667 20773
rect 263701 20745 263729 20773
rect 263763 20745 263791 20773
rect 263577 11931 263605 11959
rect 263639 11931 263667 11959
rect 263701 11931 263729 11959
rect 263763 11931 263791 11959
rect 263577 11869 263605 11897
rect 263639 11869 263667 11897
rect 263701 11869 263729 11897
rect 263763 11869 263791 11897
rect 263577 11807 263605 11835
rect 263639 11807 263667 11835
rect 263701 11807 263729 11835
rect 263763 11807 263791 11835
rect 263577 11745 263605 11773
rect 263639 11745 263667 11773
rect 263701 11745 263729 11773
rect 263763 11745 263791 11773
rect 263577 2931 263605 2959
rect 263639 2931 263667 2959
rect 263701 2931 263729 2959
rect 263763 2931 263791 2959
rect 263577 2869 263605 2897
rect 263639 2869 263667 2897
rect 263701 2869 263729 2897
rect 263763 2869 263791 2897
rect 263577 2807 263605 2835
rect 263639 2807 263667 2835
rect 263701 2807 263729 2835
rect 263763 2807 263791 2835
rect 263577 2745 263605 2773
rect 263639 2745 263667 2773
rect 263701 2745 263729 2773
rect 263763 2745 263791 2773
rect 263577 876 263605 904
rect 263639 876 263667 904
rect 263701 876 263729 904
rect 263763 876 263791 904
rect 263577 814 263605 842
rect 263639 814 263667 842
rect 263701 814 263729 842
rect 263763 814 263791 842
rect 263577 752 263605 780
rect 263639 752 263667 780
rect 263701 752 263729 780
rect 263763 752 263791 780
rect 263577 690 263605 718
rect 263639 690 263667 718
rect 263701 690 263729 718
rect 263763 690 263791 718
rect 265437 299642 265465 299670
rect 265499 299642 265527 299670
rect 265561 299642 265589 299670
rect 265623 299642 265651 299670
rect 265437 299580 265465 299608
rect 265499 299580 265527 299608
rect 265561 299580 265589 299608
rect 265623 299580 265651 299608
rect 265437 299518 265465 299546
rect 265499 299518 265527 299546
rect 265561 299518 265589 299546
rect 265623 299518 265651 299546
rect 265437 299456 265465 299484
rect 265499 299456 265527 299484
rect 265561 299456 265589 299484
rect 265623 299456 265651 299484
rect 265437 293931 265465 293959
rect 265499 293931 265527 293959
rect 265561 293931 265589 293959
rect 265623 293931 265651 293959
rect 265437 293869 265465 293897
rect 265499 293869 265527 293897
rect 265561 293869 265589 293897
rect 265623 293869 265651 293897
rect 265437 293807 265465 293835
rect 265499 293807 265527 293835
rect 265561 293807 265589 293835
rect 265623 293807 265651 293835
rect 265437 293745 265465 293773
rect 265499 293745 265527 293773
rect 265561 293745 265589 293773
rect 265623 293745 265651 293773
rect 265437 284931 265465 284959
rect 265499 284931 265527 284959
rect 265561 284931 265589 284959
rect 265623 284931 265651 284959
rect 265437 284869 265465 284897
rect 265499 284869 265527 284897
rect 265561 284869 265589 284897
rect 265623 284869 265651 284897
rect 265437 284807 265465 284835
rect 265499 284807 265527 284835
rect 265561 284807 265589 284835
rect 265623 284807 265651 284835
rect 265437 284745 265465 284773
rect 265499 284745 265527 284773
rect 265561 284745 265589 284773
rect 265623 284745 265651 284773
rect 265437 275931 265465 275959
rect 265499 275931 265527 275959
rect 265561 275931 265589 275959
rect 265623 275931 265651 275959
rect 265437 275869 265465 275897
rect 265499 275869 265527 275897
rect 265561 275869 265589 275897
rect 265623 275869 265651 275897
rect 265437 275807 265465 275835
rect 265499 275807 265527 275835
rect 265561 275807 265589 275835
rect 265623 275807 265651 275835
rect 265437 275745 265465 275773
rect 265499 275745 265527 275773
rect 265561 275745 265589 275773
rect 265623 275745 265651 275773
rect 265437 266931 265465 266959
rect 265499 266931 265527 266959
rect 265561 266931 265589 266959
rect 265623 266931 265651 266959
rect 265437 266869 265465 266897
rect 265499 266869 265527 266897
rect 265561 266869 265589 266897
rect 265623 266869 265651 266897
rect 265437 266807 265465 266835
rect 265499 266807 265527 266835
rect 265561 266807 265589 266835
rect 265623 266807 265651 266835
rect 265437 266745 265465 266773
rect 265499 266745 265527 266773
rect 265561 266745 265589 266773
rect 265623 266745 265651 266773
rect 265437 257931 265465 257959
rect 265499 257931 265527 257959
rect 265561 257931 265589 257959
rect 265623 257931 265651 257959
rect 265437 257869 265465 257897
rect 265499 257869 265527 257897
rect 265561 257869 265589 257897
rect 265623 257869 265651 257897
rect 265437 257807 265465 257835
rect 265499 257807 265527 257835
rect 265561 257807 265589 257835
rect 265623 257807 265651 257835
rect 265437 257745 265465 257773
rect 265499 257745 265527 257773
rect 265561 257745 265589 257773
rect 265623 257745 265651 257773
rect 265437 248931 265465 248959
rect 265499 248931 265527 248959
rect 265561 248931 265589 248959
rect 265623 248931 265651 248959
rect 265437 248869 265465 248897
rect 265499 248869 265527 248897
rect 265561 248869 265589 248897
rect 265623 248869 265651 248897
rect 265437 248807 265465 248835
rect 265499 248807 265527 248835
rect 265561 248807 265589 248835
rect 265623 248807 265651 248835
rect 265437 248745 265465 248773
rect 265499 248745 265527 248773
rect 265561 248745 265589 248773
rect 265623 248745 265651 248773
rect 265437 239931 265465 239959
rect 265499 239931 265527 239959
rect 265561 239931 265589 239959
rect 265623 239931 265651 239959
rect 265437 239869 265465 239897
rect 265499 239869 265527 239897
rect 265561 239869 265589 239897
rect 265623 239869 265651 239897
rect 265437 239807 265465 239835
rect 265499 239807 265527 239835
rect 265561 239807 265589 239835
rect 265623 239807 265651 239835
rect 265437 239745 265465 239773
rect 265499 239745 265527 239773
rect 265561 239745 265589 239773
rect 265623 239745 265651 239773
rect 265437 230931 265465 230959
rect 265499 230931 265527 230959
rect 265561 230931 265589 230959
rect 265623 230931 265651 230959
rect 265437 230869 265465 230897
rect 265499 230869 265527 230897
rect 265561 230869 265589 230897
rect 265623 230869 265651 230897
rect 265437 230807 265465 230835
rect 265499 230807 265527 230835
rect 265561 230807 265589 230835
rect 265623 230807 265651 230835
rect 265437 230745 265465 230773
rect 265499 230745 265527 230773
rect 265561 230745 265589 230773
rect 265623 230745 265651 230773
rect 265437 221931 265465 221959
rect 265499 221931 265527 221959
rect 265561 221931 265589 221959
rect 265623 221931 265651 221959
rect 265437 221869 265465 221897
rect 265499 221869 265527 221897
rect 265561 221869 265589 221897
rect 265623 221869 265651 221897
rect 265437 221807 265465 221835
rect 265499 221807 265527 221835
rect 265561 221807 265589 221835
rect 265623 221807 265651 221835
rect 265437 221745 265465 221773
rect 265499 221745 265527 221773
rect 265561 221745 265589 221773
rect 265623 221745 265651 221773
rect 265437 212931 265465 212959
rect 265499 212931 265527 212959
rect 265561 212931 265589 212959
rect 265623 212931 265651 212959
rect 265437 212869 265465 212897
rect 265499 212869 265527 212897
rect 265561 212869 265589 212897
rect 265623 212869 265651 212897
rect 265437 212807 265465 212835
rect 265499 212807 265527 212835
rect 265561 212807 265589 212835
rect 265623 212807 265651 212835
rect 265437 212745 265465 212773
rect 265499 212745 265527 212773
rect 265561 212745 265589 212773
rect 265623 212745 265651 212773
rect 265437 203931 265465 203959
rect 265499 203931 265527 203959
rect 265561 203931 265589 203959
rect 265623 203931 265651 203959
rect 265437 203869 265465 203897
rect 265499 203869 265527 203897
rect 265561 203869 265589 203897
rect 265623 203869 265651 203897
rect 265437 203807 265465 203835
rect 265499 203807 265527 203835
rect 265561 203807 265589 203835
rect 265623 203807 265651 203835
rect 265437 203745 265465 203773
rect 265499 203745 265527 203773
rect 265561 203745 265589 203773
rect 265623 203745 265651 203773
rect 265437 194931 265465 194959
rect 265499 194931 265527 194959
rect 265561 194931 265589 194959
rect 265623 194931 265651 194959
rect 265437 194869 265465 194897
rect 265499 194869 265527 194897
rect 265561 194869 265589 194897
rect 265623 194869 265651 194897
rect 265437 194807 265465 194835
rect 265499 194807 265527 194835
rect 265561 194807 265589 194835
rect 265623 194807 265651 194835
rect 265437 194745 265465 194773
rect 265499 194745 265527 194773
rect 265561 194745 265589 194773
rect 265623 194745 265651 194773
rect 265437 185931 265465 185959
rect 265499 185931 265527 185959
rect 265561 185931 265589 185959
rect 265623 185931 265651 185959
rect 265437 185869 265465 185897
rect 265499 185869 265527 185897
rect 265561 185869 265589 185897
rect 265623 185869 265651 185897
rect 265437 185807 265465 185835
rect 265499 185807 265527 185835
rect 265561 185807 265589 185835
rect 265623 185807 265651 185835
rect 265437 185745 265465 185773
rect 265499 185745 265527 185773
rect 265561 185745 265589 185773
rect 265623 185745 265651 185773
rect 265437 176931 265465 176959
rect 265499 176931 265527 176959
rect 265561 176931 265589 176959
rect 265623 176931 265651 176959
rect 265437 176869 265465 176897
rect 265499 176869 265527 176897
rect 265561 176869 265589 176897
rect 265623 176869 265651 176897
rect 265437 176807 265465 176835
rect 265499 176807 265527 176835
rect 265561 176807 265589 176835
rect 265623 176807 265651 176835
rect 265437 176745 265465 176773
rect 265499 176745 265527 176773
rect 265561 176745 265589 176773
rect 265623 176745 265651 176773
rect 265437 167931 265465 167959
rect 265499 167931 265527 167959
rect 265561 167931 265589 167959
rect 265623 167931 265651 167959
rect 265437 167869 265465 167897
rect 265499 167869 265527 167897
rect 265561 167869 265589 167897
rect 265623 167869 265651 167897
rect 265437 167807 265465 167835
rect 265499 167807 265527 167835
rect 265561 167807 265589 167835
rect 265623 167807 265651 167835
rect 265437 167745 265465 167773
rect 265499 167745 265527 167773
rect 265561 167745 265589 167773
rect 265623 167745 265651 167773
rect 265437 158931 265465 158959
rect 265499 158931 265527 158959
rect 265561 158931 265589 158959
rect 265623 158931 265651 158959
rect 265437 158869 265465 158897
rect 265499 158869 265527 158897
rect 265561 158869 265589 158897
rect 265623 158869 265651 158897
rect 265437 158807 265465 158835
rect 265499 158807 265527 158835
rect 265561 158807 265589 158835
rect 265623 158807 265651 158835
rect 265437 158745 265465 158773
rect 265499 158745 265527 158773
rect 265561 158745 265589 158773
rect 265623 158745 265651 158773
rect 265437 149931 265465 149959
rect 265499 149931 265527 149959
rect 265561 149931 265589 149959
rect 265623 149931 265651 149959
rect 265437 149869 265465 149897
rect 265499 149869 265527 149897
rect 265561 149869 265589 149897
rect 265623 149869 265651 149897
rect 265437 149807 265465 149835
rect 265499 149807 265527 149835
rect 265561 149807 265589 149835
rect 265623 149807 265651 149835
rect 265437 149745 265465 149773
rect 265499 149745 265527 149773
rect 265561 149745 265589 149773
rect 265623 149745 265651 149773
rect 265437 140931 265465 140959
rect 265499 140931 265527 140959
rect 265561 140931 265589 140959
rect 265623 140931 265651 140959
rect 265437 140869 265465 140897
rect 265499 140869 265527 140897
rect 265561 140869 265589 140897
rect 265623 140869 265651 140897
rect 265437 140807 265465 140835
rect 265499 140807 265527 140835
rect 265561 140807 265589 140835
rect 265623 140807 265651 140835
rect 265437 140745 265465 140773
rect 265499 140745 265527 140773
rect 265561 140745 265589 140773
rect 265623 140745 265651 140773
rect 265437 131931 265465 131959
rect 265499 131931 265527 131959
rect 265561 131931 265589 131959
rect 265623 131931 265651 131959
rect 265437 131869 265465 131897
rect 265499 131869 265527 131897
rect 265561 131869 265589 131897
rect 265623 131869 265651 131897
rect 265437 131807 265465 131835
rect 265499 131807 265527 131835
rect 265561 131807 265589 131835
rect 265623 131807 265651 131835
rect 265437 131745 265465 131773
rect 265499 131745 265527 131773
rect 265561 131745 265589 131773
rect 265623 131745 265651 131773
rect 265437 122931 265465 122959
rect 265499 122931 265527 122959
rect 265561 122931 265589 122959
rect 265623 122931 265651 122959
rect 265437 122869 265465 122897
rect 265499 122869 265527 122897
rect 265561 122869 265589 122897
rect 265623 122869 265651 122897
rect 265437 122807 265465 122835
rect 265499 122807 265527 122835
rect 265561 122807 265589 122835
rect 265623 122807 265651 122835
rect 265437 122745 265465 122773
rect 265499 122745 265527 122773
rect 265561 122745 265589 122773
rect 265623 122745 265651 122773
rect 265437 113931 265465 113959
rect 265499 113931 265527 113959
rect 265561 113931 265589 113959
rect 265623 113931 265651 113959
rect 265437 113869 265465 113897
rect 265499 113869 265527 113897
rect 265561 113869 265589 113897
rect 265623 113869 265651 113897
rect 265437 113807 265465 113835
rect 265499 113807 265527 113835
rect 265561 113807 265589 113835
rect 265623 113807 265651 113835
rect 265437 113745 265465 113773
rect 265499 113745 265527 113773
rect 265561 113745 265589 113773
rect 265623 113745 265651 113773
rect 265437 104931 265465 104959
rect 265499 104931 265527 104959
rect 265561 104931 265589 104959
rect 265623 104931 265651 104959
rect 265437 104869 265465 104897
rect 265499 104869 265527 104897
rect 265561 104869 265589 104897
rect 265623 104869 265651 104897
rect 265437 104807 265465 104835
rect 265499 104807 265527 104835
rect 265561 104807 265589 104835
rect 265623 104807 265651 104835
rect 265437 104745 265465 104773
rect 265499 104745 265527 104773
rect 265561 104745 265589 104773
rect 265623 104745 265651 104773
rect 265437 95931 265465 95959
rect 265499 95931 265527 95959
rect 265561 95931 265589 95959
rect 265623 95931 265651 95959
rect 265437 95869 265465 95897
rect 265499 95869 265527 95897
rect 265561 95869 265589 95897
rect 265623 95869 265651 95897
rect 265437 95807 265465 95835
rect 265499 95807 265527 95835
rect 265561 95807 265589 95835
rect 265623 95807 265651 95835
rect 265437 95745 265465 95773
rect 265499 95745 265527 95773
rect 265561 95745 265589 95773
rect 265623 95745 265651 95773
rect 265437 86931 265465 86959
rect 265499 86931 265527 86959
rect 265561 86931 265589 86959
rect 265623 86931 265651 86959
rect 265437 86869 265465 86897
rect 265499 86869 265527 86897
rect 265561 86869 265589 86897
rect 265623 86869 265651 86897
rect 265437 86807 265465 86835
rect 265499 86807 265527 86835
rect 265561 86807 265589 86835
rect 265623 86807 265651 86835
rect 265437 86745 265465 86773
rect 265499 86745 265527 86773
rect 265561 86745 265589 86773
rect 265623 86745 265651 86773
rect 265437 77931 265465 77959
rect 265499 77931 265527 77959
rect 265561 77931 265589 77959
rect 265623 77931 265651 77959
rect 265437 77869 265465 77897
rect 265499 77869 265527 77897
rect 265561 77869 265589 77897
rect 265623 77869 265651 77897
rect 265437 77807 265465 77835
rect 265499 77807 265527 77835
rect 265561 77807 265589 77835
rect 265623 77807 265651 77835
rect 265437 77745 265465 77773
rect 265499 77745 265527 77773
rect 265561 77745 265589 77773
rect 265623 77745 265651 77773
rect 265437 68931 265465 68959
rect 265499 68931 265527 68959
rect 265561 68931 265589 68959
rect 265623 68931 265651 68959
rect 265437 68869 265465 68897
rect 265499 68869 265527 68897
rect 265561 68869 265589 68897
rect 265623 68869 265651 68897
rect 265437 68807 265465 68835
rect 265499 68807 265527 68835
rect 265561 68807 265589 68835
rect 265623 68807 265651 68835
rect 265437 68745 265465 68773
rect 265499 68745 265527 68773
rect 265561 68745 265589 68773
rect 265623 68745 265651 68773
rect 265437 59931 265465 59959
rect 265499 59931 265527 59959
rect 265561 59931 265589 59959
rect 265623 59931 265651 59959
rect 265437 59869 265465 59897
rect 265499 59869 265527 59897
rect 265561 59869 265589 59897
rect 265623 59869 265651 59897
rect 265437 59807 265465 59835
rect 265499 59807 265527 59835
rect 265561 59807 265589 59835
rect 265623 59807 265651 59835
rect 265437 59745 265465 59773
rect 265499 59745 265527 59773
rect 265561 59745 265589 59773
rect 265623 59745 265651 59773
rect 265437 50931 265465 50959
rect 265499 50931 265527 50959
rect 265561 50931 265589 50959
rect 265623 50931 265651 50959
rect 265437 50869 265465 50897
rect 265499 50869 265527 50897
rect 265561 50869 265589 50897
rect 265623 50869 265651 50897
rect 265437 50807 265465 50835
rect 265499 50807 265527 50835
rect 265561 50807 265589 50835
rect 265623 50807 265651 50835
rect 265437 50745 265465 50773
rect 265499 50745 265527 50773
rect 265561 50745 265589 50773
rect 265623 50745 265651 50773
rect 265437 41931 265465 41959
rect 265499 41931 265527 41959
rect 265561 41931 265589 41959
rect 265623 41931 265651 41959
rect 265437 41869 265465 41897
rect 265499 41869 265527 41897
rect 265561 41869 265589 41897
rect 265623 41869 265651 41897
rect 265437 41807 265465 41835
rect 265499 41807 265527 41835
rect 265561 41807 265589 41835
rect 265623 41807 265651 41835
rect 265437 41745 265465 41773
rect 265499 41745 265527 41773
rect 265561 41745 265589 41773
rect 265623 41745 265651 41773
rect 265437 32931 265465 32959
rect 265499 32931 265527 32959
rect 265561 32931 265589 32959
rect 265623 32931 265651 32959
rect 265437 32869 265465 32897
rect 265499 32869 265527 32897
rect 265561 32869 265589 32897
rect 265623 32869 265651 32897
rect 265437 32807 265465 32835
rect 265499 32807 265527 32835
rect 265561 32807 265589 32835
rect 265623 32807 265651 32835
rect 265437 32745 265465 32773
rect 265499 32745 265527 32773
rect 265561 32745 265589 32773
rect 265623 32745 265651 32773
rect 265437 23931 265465 23959
rect 265499 23931 265527 23959
rect 265561 23931 265589 23959
rect 265623 23931 265651 23959
rect 265437 23869 265465 23897
rect 265499 23869 265527 23897
rect 265561 23869 265589 23897
rect 265623 23869 265651 23897
rect 265437 23807 265465 23835
rect 265499 23807 265527 23835
rect 265561 23807 265589 23835
rect 265623 23807 265651 23835
rect 265437 23745 265465 23773
rect 265499 23745 265527 23773
rect 265561 23745 265589 23773
rect 265623 23745 265651 23773
rect 265437 14931 265465 14959
rect 265499 14931 265527 14959
rect 265561 14931 265589 14959
rect 265623 14931 265651 14959
rect 265437 14869 265465 14897
rect 265499 14869 265527 14897
rect 265561 14869 265589 14897
rect 265623 14869 265651 14897
rect 265437 14807 265465 14835
rect 265499 14807 265527 14835
rect 265561 14807 265589 14835
rect 265623 14807 265651 14835
rect 265437 14745 265465 14773
rect 265499 14745 265527 14773
rect 265561 14745 265589 14773
rect 265623 14745 265651 14773
rect 265437 5931 265465 5959
rect 265499 5931 265527 5959
rect 265561 5931 265589 5959
rect 265623 5931 265651 5959
rect 265437 5869 265465 5897
rect 265499 5869 265527 5897
rect 265561 5869 265589 5897
rect 265623 5869 265651 5897
rect 265437 5807 265465 5835
rect 265499 5807 265527 5835
rect 265561 5807 265589 5835
rect 265623 5807 265651 5835
rect 265437 5745 265465 5773
rect 265499 5745 265527 5773
rect 265561 5745 265589 5773
rect 265623 5745 265651 5773
rect 265437 396 265465 424
rect 265499 396 265527 424
rect 265561 396 265589 424
rect 265623 396 265651 424
rect 265437 334 265465 362
rect 265499 334 265527 362
rect 265561 334 265589 362
rect 265623 334 265651 362
rect 265437 272 265465 300
rect 265499 272 265527 300
rect 265561 272 265589 300
rect 265623 272 265651 300
rect 265437 210 265465 238
rect 265499 210 265527 238
rect 265561 210 265589 238
rect 265623 210 265651 238
rect 272577 299162 272605 299190
rect 272639 299162 272667 299190
rect 272701 299162 272729 299190
rect 272763 299162 272791 299190
rect 272577 299100 272605 299128
rect 272639 299100 272667 299128
rect 272701 299100 272729 299128
rect 272763 299100 272791 299128
rect 272577 299038 272605 299066
rect 272639 299038 272667 299066
rect 272701 299038 272729 299066
rect 272763 299038 272791 299066
rect 272577 298976 272605 299004
rect 272639 298976 272667 299004
rect 272701 298976 272729 299004
rect 272763 298976 272791 299004
rect 272577 290931 272605 290959
rect 272639 290931 272667 290959
rect 272701 290931 272729 290959
rect 272763 290931 272791 290959
rect 272577 290869 272605 290897
rect 272639 290869 272667 290897
rect 272701 290869 272729 290897
rect 272763 290869 272791 290897
rect 272577 290807 272605 290835
rect 272639 290807 272667 290835
rect 272701 290807 272729 290835
rect 272763 290807 272791 290835
rect 272577 290745 272605 290773
rect 272639 290745 272667 290773
rect 272701 290745 272729 290773
rect 272763 290745 272791 290773
rect 272577 281931 272605 281959
rect 272639 281931 272667 281959
rect 272701 281931 272729 281959
rect 272763 281931 272791 281959
rect 272577 281869 272605 281897
rect 272639 281869 272667 281897
rect 272701 281869 272729 281897
rect 272763 281869 272791 281897
rect 272577 281807 272605 281835
rect 272639 281807 272667 281835
rect 272701 281807 272729 281835
rect 272763 281807 272791 281835
rect 272577 281745 272605 281773
rect 272639 281745 272667 281773
rect 272701 281745 272729 281773
rect 272763 281745 272791 281773
rect 272577 272931 272605 272959
rect 272639 272931 272667 272959
rect 272701 272931 272729 272959
rect 272763 272931 272791 272959
rect 272577 272869 272605 272897
rect 272639 272869 272667 272897
rect 272701 272869 272729 272897
rect 272763 272869 272791 272897
rect 272577 272807 272605 272835
rect 272639 272807 272667 272835
rect 272701 272807 272729 272835
rect 272763 272807 272791 272835
rect 272577 272745 272605 272773
rect 272639 272745 272667 272773
rect 272701 272745 272729 272773
rect 272763 272745 272791 272773
rect 272577 263931 272605 263959
rect 272639 263931 272667 263959
rect 272701 263931 272729 263959
rect 272763 263931 272791 263959
rect 272577 263869 272605 263897
rect 272639 263869 272667 263897
rect 272701 263869 272729 263897
rect 272763 263869 272791 263897
rect 272577 263807 272605 263835
rect 272639 263807 272667 263835
rect 272701 263807 272729 263835
rect 272763 263807 272791 263835
rect 272577 263745 272605 263773
rect 272639 263745 272667 263773
rect 272701 263745 272729 263773
rect 272763 263745 272791 263773
rect 272577 254931 272605 254959
rect 272639 254931 272667 254959
rect 272701 254931 272729 254959
rect 272763 254931 272791 254959
rect 272577 254869 272605 254897
rect 272639 254869 272667 254897
rect 272701 254869 272729 254897
rect 272763 254869 272791 254897
rect 272577 254807 272605 254835
rect 272639 254807 272667 254835
rect 272701 254807 272729 254835
rect 272763 254807 272791 254835
rect 272577 254745 272605 254773
rect 272639 254745 272667 254773
rect 272701 254745 272729 254773
rect 272763 254745 272791 254773
rect 272577 245931 272605 245959
rect 272639 245931 272667 245959
rect 272701 245931 272729 245959
rect 272763 245931 272791 245959
rect 272577 245869 272605 245897
rect 272639 245869 272667 245897
rect 272701 245869 272729 245897
rect 272763 245869 272791 245897
rect 272577 245807 272605 245835
rect 272639 245807 272667 245835
rect 272701 245807 272729 245835
rect 272763 245807 272791 245835
rect 272577 245745 272605 245773
rect 272639 245745 272667 245773
rect 272701 245745 272729 245773
rect 272763 245745 272791 245773
rect 272577 236931 272605 236959
rect 272639 236931 272667 236959
rect 272701 236931 272729 236959
rect 272763 236931 272791 236959
rect 272577 236869 272605 236897
rect 272639 236869 272667 236897
rect 272701 236869 272729 236897
rect 272763 236869 272791 236897
rect 272577 236807 272605 236835
rect 272639 236807 272667 236835
rect 272701 236807 272729 236835
rect 272763 236807 272791 236835
rect 272577 236745 272605 236773
rect 272639 236745 272667 236773
rect 272701 236745 272729 236773
rect 272763 236745 272791 236773
rect 272577 227931 272605 227959
rect 272639 227931 272667 227959
rect 272701 227931 272729 227959
rect 272763 227931 272791 227959
rect 272577 227869 272605 227897
rect 272639 227869 272667 227897
rect 272701 227869 272729 227897
rect 272763 227869 272791 227897
rect 272577 227807 272605 227835
rect 272639 227807 272667 227835
rect 272701 227807 272729 227835
rect 272763 227807 272791 227835
rect 272577 227745 272605 227773
rect 272639 227745 272667 227773
rect 272701 227745 272729 227773
rect 272763 227745 272791 227773
rect 272577 218931 272605 218959
rect 272639 218931 272667 218959
rect 272701 218931 272729 218959
rect 272763 218931 272791 218959
rect 272577 218869 272605 218897
rect 272639 218869 272667 218897
rect 272701 218869 272729 218897
rect 272763 218869 272791 218897
rect 272577 218807 272605 218835
rect 272639 218807 272667 218835
rect 272701 218807 272729 218835
rect 272763 218807 272791 218835
rect 272577 218745 272605 218773
rect 272639 218745 272667 218773
rect 272701 218745 272729 218773
rect 272763 218745 272791 218773
rect 272577 209931 272605 209959
rect 272639 209931 272667 209959
rect 272701 209931 272729 209959
rect 272763 209931 272791 209959
rect 272577 209869 272605 209897
rect 272639 209869 272667 209897
rect 272701 209869 272729 209897
rect 272763 209869 272791 209897
rect 272577 209807 272605 209835
rect 272639 209807 272667 209835
rect 272701 209807 272729 209835
rect 272763 209807 272791 209835
rect 272577 209745 272605 209773
rect 272639 209745 272667 209773
rect 272701 209745 272729 209773
rect 272763 209745 272791 209773
rect 272577 200931 272605 200959
rect 272639 200931 272667 200959
rect 272701 200931 272729 200959
rect 272763 200931 272791 200959
rect 272577 200869 272605 200897
rect 272639 200869 272667 200897
rect 272701 200869 272729 200897
rect 272763 200869 272791 200897
rect 272577 200807 272605 200835
rect 272639 200807 272667 200835
rect 272701 200807 272729 200835
rect 272763 200807 272791 200835
rect 272577 200745 272605 200773
rect 272639 200745 272667 200773
rect 272701 200745 272729 200773
rect 272763 200745 272791 200773
rect 272577 191931 272605 191959
rect 272639 191931 272667 191959
rect 272701 191931 272729 191959
rect 272763 191931 272791 191959
rect 272577 191869 272605 191897
rect 272639 191869 272667 191897
rect 272701 191869 272729 191897
rect 272763 191869 272791 191897
rect 272577 191807 272605 191835
rect 272639 191807 272667 191835
rect 272701 191807 272729 191835
rect 272763 191807 272791 191835
rect 272577 191745 272605 191773
rect 272639 191745 272667 191773
rect 272701 191745 272729 191773
rect 272763 191745 272791 191773
rect 272577 182931 272605 182959
rect 272639 182931 272667 182959
rect 272701 182931 272729 182959
rect 272763 182931 272791 182959
rect 272577 182869 272605 182897
rect 272639 182869 272667 182897
rect 272701 182869 272729 182897
rect 272763 182869 272791 182897
rect 272577 182807 272605 182835
rect 272639 182807 272667 182835
rect 272701 182807 272729 182835
rect 272763 182807 272791 182835
rect 272577 182745 272605 182773
rect 272639 182745 272667 182773
rect 272701 182745 272729 182773
rect 272763 182745 272791 182773
rect 272577 173931 272605 173959
rect 272639 173931 272667 173959
rect 272701 173931 272729 173959
rect 272763 173931 272791 173959
rect 272577 173869 272605 173897
rect 272639 173869 272667 173897
rect 272701 173869 272729 173897
rect 272763 173869 272791 173897
rect 272577 173807 272605 173835
rect 272639 173807 272667 173835
rect 272701 173807 272729 173835
rect 272763 173807 272791 173835
rect 272577 173745 272605 173773
rect 272639 173745 272667 173773
rect 272701 173745 272729 173773
rect 272763 173745 272791 173773
rect 272577 164931 272605 164959
rect 272639 164931 272667 164959
rect 272701 164931 272729 164959
rect 272763 164931 272791 164959
rect 272577 164869 272605 164897
rect 272639 164869 272667 164897
rect 272701 164869 272729 164897
rect 272763 164869 272791 164897
rect 272577 164807 272605 164835
rect 272639 164807 272667 164835
rect 272701 164807 272729 164835
rect 272763 164807 272791 164835
rect 272577 164745 272605 164773
rect 272639 164745 272667 164773
rect 272701 164745 272729 164773
rect 272763 164745 272791 164773
rect 272577 155931 272605 155959
rect 272639 155931 272667 155959
rect 272701 155931 272729 155959
rect 272763 155931 272791 155959
rect 272577 155869 272605 155897
rect 272639 155869 272667 155897
rect 272701 155869 272729 155897
rect 272763 155869 272791 155897
rect 272577 155807 272605 155835
rect 272639 155807 272667 155835
rect 272701 155807 272729 155835
rect 272763 155807 272791 155835
rect 272577 155745 272605 155773
rect 272639 155745 272667 155773
rect 272701 155745 272729 155773
rect 272763 155745 272791 155773
rect 272577 146931 272605 146959
rect 272639 146931 272667 146959
rect 272701 146931 272729 146959
rect 272763 146931 272791 146959
rect 272577 146869 272605 146897
rect 272639 146869 272667 146897
rect 272701 146869 272729 146897
rect 272763 146869 272791 146897
rect 272577 146807 272605 146835
rect 272639 146807 272667 146835
rect 272701 146807 272729 146835
rect 272763 146807 272791 146835
rect 272577 146745 272605 146773
rect 272639 146745 272667 146773
rect 272701 146745 272729 146773
rect 272763 146745 272791 146773
rect 272577 137931 272605 137959
rect 272639 137931 272667 137959
rect 272701 137931 272729 137959
rect 272763 137931 272791 137959
rect 272577 137869 272605 137897
rect 272639 137869 272667 137897
rect 272701 137869 272729 137897
rect 272763 137869 272791 137897
rect 272577 137807 272605 137835
rect 272639 137807 272667 137835
rect 272701 137807 272729 137835
rect 272763 137807 272791 137835
rect 272577 137745 272605 137773
rect 272639 137745 272667 137773
rect 272701 137745 272729 137773
rect 272763 137745 272791 137773
rect 272577 128931 272605 128959
rect 272639 128931 272667 128959
rect 272701 128931 272729 128959
rect 272763 128931 272791 128959
rect 272577 128869 272605 128897
rect 272639 128869 272667 128897
rect 272701 128869 272729 128897
rect 272763 128869 272791 128897
rect 272577 128807 272605 128835
rect 272639 128807 272667 128835
rect 272701 128807 272729 128835
rect 272763 128807 272791 128835
rect 272577 128745 272605 128773
rect 272639 128745 272667 128773
rect 272701 128745 272729 128773
rect 272763 128745 272791 128773
rect 272577 119931 272605 119959
rect 272639 119931 272667 119959
rect 272701 119931 272729 119959
rect 272763 119931 272791 119959
rect 272577 119869 272605 119897
rect 272639 119869 272667 119897
rect 272701 119869 272729 119897
rect 272763 119869 272791 119897
rect 272577 119807 272605 119835
rect 272639 119807 272667 119835
rect 272701 119807 272729 119835
rect 272763 119807 272791 119835
rect 272577 119745 272605 119773
rect 272639 119745 272667 119773
rect 272701 119745 272729 119773
rect 272763 119745 272791 119773
rect 272577 110931 272605 110959
rect 272639 110931 272667 110959
rect 272701 110931 272729 110959
rect 272763 110931 272791 110959
rect 272577 110869 272605 110897
rect 272639 110869 272667 110897
rect 272701 110869 272729 110897
rect 272763 110869 272791 110897
rect 272577 110807 272605 110835
rect 272639 110807 272667 110835
rect 272701 110807 272729 110835
rect 272763 110807 272791 110835
rect 272577 110745 272605 110773
rect 272639 110745 272667 110773
rect 272701 110745 272729 110773
rect 272763 110745 272791 110773
rect 272577 101931 272605 101959
rect 272639 101931 272667 101959
rect 272701 101931 272729 101959
rect 272763 101931 272791 101959
rect 272577 101869 272605 101897
rect 272639 101869 272667 101897
rect 272701 101869 272729 101897
rect 272763 101869 272791 101897
rect 272577 101807 272605 101835
rect 272639 101807 272667 101835
rect 272701 101807 272729 101835
rect 272763 101807 272791 101835
rect 272577 101745 272605 101773
rect 272639 101745 272667 101773
rect 272701 101745 272729 101773
rect 272763 101745 272791 101773
rect 272577 92931 272605 92959
rect 272639 92931 272667 92959
rect 272701 92931 272729 92959
rect 272763 92931 272791 92959
rect 272577 92869 272605 92897
rect 272639 92869 272667 92897
rect 272701 92869 272729 92897
rect 272763 92869 272791 92897
rect 272577 92807 272605 92835
rect 272639 92807 272667 92835
rect 272701 92807 272729 92835
rect 272763 92807 272791 92835
rect 272577 92745 272605 92773
rect 272639 92745 272667 92773
rect 272701 92745 272729 92773
rect 272763 92745 272791 92773
rect 272577 83931 272605 83959
rect 272639 83931 272667 83959
rect 272701 83931 272729 83959
rect 272763 83931 272791 83959
rect 272577 83869 272605 83897
rect 272639 83869 272667 83897
rect 272701 83869 272729 83897
rect 272763 83869 272791 83897
rect 272577 83807 272605 83835
rect 272639 83807 272667 83835
rect 272701 83807 272729 83835
rect 272763 83807 272791 83835
rect 272577 83745 272605 83773
rect 272639 83745 272667 83773
rect 272701 83745 272729 83773
rect 272763 83745 272791 83773
rect 272577 74931 272605 74959
rect 272639 74931 272667 74959
rect 272701 74931 272729 74959
rect 272763 74931 272791 74959
rect 272577 74869 272605 74897
rect 272639 74869 272667 74897
rect 272701 74869 272729 74897
rect 272763 74869 272791 74897
rect 272577 74807 272605 74835
rect 272639 74807 272667 74835
rect 272701 74807 272729 74835
rect 272763 74807 272791 74835
rect 272577 74745 272605 74773
rect 272639 74745 272667 74773
rect 272701 74745 272729 74773
rect 272763 74745 272791 74773
rect 272577 65931 272605 65959
rect 272639 65931 272667 65959
rect 272701 65931 272729 65959
rect 272763 65931 272791 65959
rect 272577 65869 272605 65897
rect 272639 65869 272667 65897
rect 272701 65869 272729 65897
rect 272763 65869 272791 65897
rect 272577 65807 272605 65835
rect 272639 65807 272667 65835
rect 272701 65807 272729 65835
rect 272763 65807 272791 65835
rect 272577 65745 272605 65773
rect 272639 65745 272667 65773
rect 272701 65745 272729 65773
rect 272763 65745 272791 65773
rect 272577 56931 272605 56959
rect 272639 56931 272667 56959
rect 272701 56931 272729 56959
rect 272763 56931 272791 56959
rect 272577 56869 272605 56897
rect 272639 56869 272667 56897
rect 272701 56869 272729 56897
rect 272763 56869 272791 56897
rect 272577 56807 272605 56835
rect 272639 56807 272667 56835
rect 272701 56807 272729 56835
rect 272763 56807 272791 56835
rect 272577 56745 272605 56773
rect 272639 56745 272667 56773
rect 272701 56745 272729 56773
rect 272763 56745 272791 56773
rect 272577 47931 272605 47959
rect 272639 47931 272667 47959
rect 272701 47931 272729 47959
rect 272763 47931 272791 47959
rect 272577 47869 272605 47897
rect 272639 47869 272667 47897
rect 272701 47869 272729 47897
rect 272763 47869 272791 47897
rect 272577 47807 272605 47835
rect 272639 47807 272667 47835
rect 272701 47807 272729 47835
rect 272763 47807 272791 47835
rect 272577 47745 272605 47773
rect 272639 47745 272667 47773
rect 272701 47745 272729 47773
rect 272763 47745 272791 47773
rect 272577 38931 272605 38959
rect 272639 38931 272667 38959
rect 272701 38931 272729 38959
rect 272763 38931 272791 38959
rect 272577 38869 272605 38897
rect 272639 38869 272667 38897
rect 272701 38869 272729 38897
rect 272763 38869 272791 38897
rect 272577 38807 272605 38835
rect 272639 38807 272667 38835
rect 272701 38807 272729 38835
rect 272763 38807 272791 38835
rect 272577 38745 272605 38773
rect 272639 38745 272667 38773
rect 272701 38745 272729 38773
rect 272763 38745 272791 38773
rect 272577 29931 272605 29959
rect 272639 29931 272667 29959
rect 272701 29931 272729 29959
rect 272763 29931 272791 29959
rect 272577 29869 272605 29897
rect 272639 29869 272667 29897
rect 272701 29869 272729 29897
rect 272763 29869 272791 29897
rect 272577 29807 272605 29835
rect 272639 29807 272667 29835
rect 272701 29807 272729 29835
rect 272763 29807 272791 29835
rect 272577 29745 272605 29773
rect 272639 29745 272667 29773
rect 272701 29745 272729 29773
rect 272763 29745 272791 29773
rect 272577 20931 272605 20959
rect 272639 20931 272667 20959
rect 272701 20931 272729 20959
rect 272763 20931 272791 20959
rect 272577 20869 272605 20897
rect 272639 20869 272667 20897
rect 272701 20869 272729 20897
rect 272763 20869 272791 20897
rect 272577 20807 272605 20835
rect 272639 20807 272667 20835
rect 272701 20807 272729 20835
rect 272763 20807 272791 20835
rect 272577 20745 272605 20773
rect 272639 20745 272667 20773
rect 272701 20745 272729 20773
rect 272763 20745 272791 20773
rect 272577 11931 272605 11959
rect 272639 11931 272667 11959
rect 272701 11931 272729 11959
rect 272763 11931 272791 11959
rect 272577 11869 272605 11897
rect 272639 11869 272667 11897
rect 272701 11869 272729 11897
rect 272763 11869 272791 11897
rect 272577 11807 272605 11835
rect 272639 11807 272667 11835
rect 272701 11807 272729 11835
rect 272763 11807 272791 11835
rect 272577 11745 272605 11773
rect 272639 11745 272667 11773
rect 272701 11745 272729 11773
rect 272763 11745 272791 11773
rect 272577 2931 272605 2959
rect 272639 2931 272667 2959
rect 272701 2931 272729 2959
rect 272763 2931 272791 2959
rect 272577 2869 272605 2897
rect 272639 2869 272667 2897
rect 272701 2869 272729 2897
rect 272763 2869 272791 2897
rect 272577 2807 272605 2835
rect 272639 2807 272667 2835
rect 272701 2807 272729 2835
rect 272763 2807 272791 2835
rect 272577 2745 272605 2773
rect 272639 2745 272667 2773
rect 272701 2745 272729 2773
rect 272763 2745 272791 2773
rect 272577 876 272605 904
rect 272639 876 272667 904
rect 272701 876 272729 904
rect 272763 876 272791 904
rect 272577 814 272605 842
rect 272639 814 272667 842
rect 272701 814 272729 842
rect 272763 814 272791 842
rect 272577 752 272605 780
rect 272639 752 272667 780
rect 272701 752 272729 780
rect 272763 752 272791 780
rect 272577 690 272605 718
rect 272639 690 272667 718
rect 272701 690 272729 718
rect 272763 690 272791 718
rect 274437 299642 274465 299670
rect 274499 299642 274527 299670
rect 274561 299642 274589 299670
rect 274623 299642 274651 299670
rect 274437 299580 274465 299608
rect 274499 299580 274527 299608
rect 274561 299580 274589 299608
rect 274623 299580 274651 299608
rect 274437 299518 274465 299546
rect 274499 299518 274527 299546
rect 274561 299518 274589 299546
rect 274623 299518 274651 299546
rect 274437 299456 274465 299484
rect 274499 299456 274527 299484
rect 274561 299456 274589 299484
rect 274623 299456 274651 299484
rect 274437 293931 274465 293959
rect 274499 293931 274527 293959
rect 274561 293931 274589 293959
rect 274623 293931 274651 293959
rect 274437 293869 274465 293897
rect 274499 293869 274527 293897
rect 274561 293869 274589 293897
rect 274623 293869 274651 293897
rect 274437 293807 274465 293835
rect 274499 293807 274527 293835
rect 274561 293807 274589 293835
rect 274623 293807 274651 293835
rect 274437 293745 274465 293773
rect 274499 293745 274527 293773
rect 274561 293745 274589 293773
rect 274623 293745 274651 293773
rect 274437 284931 274465 284959
rect 274499 284931 274527 284959
rect 274561 284931 274589 284959
rect 274623 284931 274651 284959
rect 274437 284869 274465 284897
rect 274499 284869 274527 284897
rect 274561 284869 274589 284897
rect 274623 284869 274651 284897
rect 274437 284807 274465 284835
rect 274499 284807 274527 284835
rect 274561 284807 274589 284835
rect 274623 284807 274651 284835
rect 274437 284745 274465 284773
rect 274499 284745 274527 284773
rect 274561 284745 274589 284773
rect 274623 284745 274651 284773
rect 274437 275931 274465 275959
rect 274499 275931 274527 275959
rect 274561 275931 274589 275959
rect 274623 275931 274651 275959
rect 274437 275869 274465 275897
rect 274499 275869 274527 275897
rect 274561 275869 274589 275897
rect 274623 275869 274651 275897
rect 274437 275807 274465 275835
rect 274499 275807 274527 275835
rect 274561 275807 274589 275835
rect 274623 275807 274651 275835
rect 274437 275745 274465 275773
rect 274499 275745 274527 275773
rect 274561 275745 274589 275773
rect 274623 275745 274651 275773
rect 274437 266931 274465 266959
rect 274499 266931 274527 266959
rect 274561 266931 274589 266959
rect 274623 266931 274651 266959
rect 274437 266869 274465 266897
rect 274499 266869 274527 266897
rect 274561 266869 274589 266897
rect 274623 266869 274651 266897
rect 274437 266807 274465 266835
rect 274499 266807 274527 266835
rect 274561 266807 274589 266835
rect 274623 266807 274651 266835
rect 274437 266745 274465 266773
rect 274499 266745 274527 266773
rect 274561 266745 274589 266773
rect 274623 266745 274651 266773
rect 274437 257931 274465 257959
rect 274499 257931 274527 257959
rect 274561 257931 274589 257959
rect 274623 257931 274651 257959
rect 274437 257869 274465 257897
rect 274499 257869 274527 257897
rect 274561 257869 274589 257897
rect 274623 257869 274651 257897
rect 274437 257807 274465 257835
rect 274499 257807 274527 257835
rect 274561 257807 274589 257835
rect 274623 257807 274651 257835
rect 274437 257745 274465 257773
rect 274499 257745 274527 257773
rect 274561 257745 274589 257773
rect 274623 257745 274651 257773
rect 274437 248931 274465 248959
rect 274499 248931 274527 248959
rect 274561 248931 274589 248959
rect 274623 248931 274651 248959
rect 274437 248869 274465 248897
rect 274499 248869 274527 248897
rect 274561 248869 274589 248897
rect 274623 248869 274651 248897
rect 274437 248807 274465 248835
rect 274499 248807 274527 248835
rect 274561 248807 274589 248835
rect 274623 248807 274651 248835
rect 274437 248745 274465 248773
rect 274499 248745 274527 248773
rect 274561 248745 274589 248773
rect 274623 248745 274651 248773
rect 274437 239931 274465 239959
rect 274499 239931 274527 239959
rect 274561 239931 274589 239959
rect 274623 239931 274651 239959
rect 274437 239869 274465 239897
rect 274499 239869 274527 239897
rect 274561 239869 274589 239897
rect 274623 239869 274651 239897
rect 274437 239807 274465 239835
rect 274499 239807 274527 239835
rect 274561 239807 274589 239835
rect 274623 239807 274651 239835
rect 274437 239745 274465 239773
rect 274499 239745 274527 239773
rect 274561 239745 274589 239773
rect 274623 239745 274651 239773
rect 274437 230931 274465 230959
rect 274499 230931 274527 230959
rect 274561 230931 274589 230959
rect 274623 230931 274651 230959
rect 274437 230869 274465 230897
rect 274499 230869 274527 230897
rect 274561 230869 274589 230897
rect 274623 230869 274651 230897
rect 274437 230807 274465 230835
rect 274499 230807 274527 230835
rect 274561 230807 274589 230835
rect 274623 230807 274651 230835
rect 274437 230745 274465 230773
rect 274499 230745 274527 230773
rect 274561 230745 274589 230773
rect 274623 230745 274651 230773
rect 274437 221931 274465 221959
rect 274499 221931 274527 221959
rect 274561 221931 274589 221959
rect 274623 221931 274651 221959
rect 274437 221869 274465 221897
rect 274499 221869 274527 221897
rect 274561 221869 274589 221897
rect 274623 221869 274651 221897
rect 274437 221807 274465 221835
rect 274499 221807 274527 221835
rect 274561 221807 274589 221835
rect 274623 221807 274651 221835
rect 274437 221745 274465 221773
rect 274499 221745 274527 221773
rect 274561 221745 274589 221773
rect 274623 221745 274651 221773
rect 274437 212931 274465 212959
rect 274499 212931 274527 212959
rect 274561 212931 274589 212959
rect 274623 212931 274651 212959
rect 274437 212869 274465 212897
rect 274499 212869 274527 212897
rect 274561 212869 274589 212897
rect 274623 212869 274651 212897
rect 274437 212807 274465 212835
rect 274499 212807 274527 212835
rect 274561 212807 274589 212835
rect 274623 212807 274651 212835
rect 274437 212745 274465 212773
rect 274499 212745 274527 212773
rect 274561 212745 274589 212773
rect 274623 212745 274651 212773
rect 274437 203931 274465 203959
rect 274499 203931 274527 203959
rect 274561 203931 274589 203959
rect 274623 203931 274651 203959
rect 274437 203869 274465 203897
rect 274499 203869 274527 203897
rect 274561 203869 274589 203897
rect 274623 203869 274651 203897
rect 274437 203807 274465 203835
rect 274499 203807 274527 203835
rect 274561 203807 274589 203835
rect 274623 203807 274651 203835
rect 274437 203745 274465 203773
rect 274499 203745 274527 203773
rect 274561 203745 274589 203773
rect 274623 203745 274651 203773
rect 274437 194931 274465 194959
rect 274499 194931 274527 194959
rect 274561 194931 274589 194959
rect 274623 194931 274651 194959
rect 274437 194869 274465 194897
rect 274499 194869 274527 194897
rect 274561 194869 274589 194897
rect 274623 194869 274651 194897
rect 274437 194807 274465 194835
rect 274499 194807 274527 194835
rect 274561 194807 274589 194835
rect 274623 194807 274651 194835
rect 274437 194745 274465 194773
rect 274499 194745 274527 194773
rect 274561 194745 274589 194773
rect 274623 194745 274651 194773
rect 274437 185931 274465 185959
rect 274499 185931 274527 185959
rect 274561 185931 274589 185959
rect 274623 185931 274651 185959
rect 274437 185869 274465 185897
rect 274499 185869 274527 185897
rect 274561 185869 274589 185897
rect 274623 185869 274651 185897
rect 274437 185807 274465 185835
rect 274499 185807 274527 185835
rect 274561 185807 274589 185835
rect 274623 185807 274651 185835
rect 274437 185745 274465 185773
rect 274499 185745 274527 185773
rect 274561 185745 274589 185773
rect 274623 185745 274651 185773
rect 274437 176931 274465 176959
rect 274499 176931 274527 176959
rect 274561 176931 274589 176959
rect 274623 176931 274651 176959
rect 274437 176869 274465 176897
rect 274499 176869 274527 176897
rect 274561 176869 274589 176897
rect 274623 176869 274651 176897
rect 274437 176807 274465 176835
rect 274499 176807 274527 176835
rect 274561 176807 274589 176835
rect 274623 176807 274651 176835
rect 274437 176745 274465 176773
rect 274499 176745 274527 176773
rect 274561 176745 274589 176773
rect 274623 176745 274651 176773
rect 274437 167931 274465 167959
rect 274499 167931 274527 167959
rect 274561 167931 274589 167959
rect 274623 167931 274651 167959
rect 274437 167869 274465 167897
rect 274499 167869 274527 167897
rect 274561 167869 274589 167897
rect 274623 167869 274651 167897
rect 274437 167807 274465 167835
rect 274499 167807 274527 167835
rect 274561 167807 274589 167835
rect 274623 167807 274651 167835
rect 274437 167745 274465 167773
rect 274499 167745 274527 167773
rect 274561 167745 274589 167773
rect 274623 167745 274651 167773
rect 274437 158931 274465 158959
rect 274499 158931 274527 158959
rect 274561 158931 274589 158959
rect 274623 158931 274651 158959
rect 274437 158869 274465 158897
rect 274499 158869 274527 158897
rect 274561 158869 274589 158897
rect 274623 158869 274651 158897
rect 274437 158807 274465 158835
rect 274499 158807 274527 158835
rect 274561 158807 274589 158835
rect 274623 158807 274651 158835
rect 274437 158745 274465 158773
rect 274499 158745 274527 158773
rect 274561 158745 274589 158773
rect 274623 158745 274651 158773
rect 274437 149931 274465 149959
rect 274499 149931 274527 149959
rect 274561 149931 274589 149959
rect 274623 149931 274651 149959
rect 274437 149869 274465 149897
rect 274499 149869 274527 149897
rect 274561 149869 274589 149897
rect 274623 149869 274651 149897
rect 274437 149807 274465 149835
rect 274499 149807 274527 149835
rect 274561 149807 274589 149835
rect 274623 149807 274651 149835
rect 274437 149745 274465 149773
rect 274499 149745 274527 149773
rect 274561 149745 274589 149773
rect 274623 149745 274651 149773
rect 274437 140931 274465 140959
rect 274499 140931 274527 140959
rect 274561 140931 274589 140959
rect 274623 140931 274651 140959
rect 274437 140869 274465 140897
rect 274499 140869 274527 140897
rect 274561 140869 274589 140897
rect 274623 140869 274651 140897
rect 274437 140807 274465 140835
rect 274499 140807 274527 140835
rect 274561 140807 274589 140835
rect 274623 140807 274651 140835
rect 274437 140745 274465 140773
rect 274499 140745 274527 140773
rect 274561 140745 274589 140773
rect 274623 140745 274651 140773
rect 274437 131931 274465 131959
rect 274499 131931 274527 131959
rect 274561 131931 274589 131959
rect 274623 131931 274651 131959
rect 274437 131869 274465 131897
rect 274499 131869 274527 131897
rect 274561 131869 274589 131897
rect 274623 131869 274651 131897
rect 274437 131807 274465 131835
rect 274499 131807 274527 131835
rect 274561 131807 274589 131835
rect 274623 131807 274651 131835
rect 274437 131745 274465 131773
rect 274499 131745 274527 131773
rect 274561 131745 274589 131773
rect 274623 131745 274651 131773
rect 274437 122931 274465 122959
rect 274499 122931 274527 122959
rect 274561 122931 274589 122959
rect 274623 122931 274651 122959
rect 274437 122869 274465 122897
rect 274499 122869 274527 122897
rect 274561 122869 274589 122897
rect 274623 122869 274651 122897
rect 274437 122807 274465 122835
rect 274499 122807 274527 122835
rect 274561 122807 274589 122835
rect 274623 122807 274651 122835
rect 274437 122745 274465 122773
rect 274499 122745 274527 122773
rect 274561 122745 274589 122773
rect 274623 122745 274651 122773
rect 274437 113931 274465 113959
rect 274499 113931 274527 113959
rect 274561 113931 274589 113959
rect 274623 113931 274651 113959
rect 274437 113869 274465 113897
rect 274499 113869 274527 113897
rect 274561 113869 274589 113897
rect 274623 113869 274651 113897
rect 274437 113807 274465 113835
rect 274499 113807 274527 113835
rect 274561 113807 274589 113835
rect 274623 113807 274651 113835
rect 274437 113745 274465 113773
rect 274499 113745 274527 113773
rect 274561 113745 274589 113773
rect 274623 113745 274651 113773
rect 274437 104931 274465 104959
rect 274499 104931 274527 104959
rect 274561 104931 274589 104959
rect 274623 104931 274651 104959
rect 274437 104869 274465 104897
rect 274499 104869 274527 104897
rect 274561 104869 274589 104897
rect 274623 104869 274651 104897
rect 274437 104807 274465 104835
rect 274499 104807 274527 104835
rect 274561 104807 274589 104835
rect 274623 104807 274651 104835
rect 274437 104745 274465 104773
rect 274499 104745 274527 104773
rect 274561 104745 274589 104773
rect 274623 104745 274651 104773
rect 274437 95931 274465 95959
rect 274499 95931 274527 95959
rect 274561 95931 274589 95959
rect 274623 95931 274651 95959
rect 274437 95869 274465 95897
rect 274499 95869 274527 95897
rect 274561 95869 274589 95897
rect 274623 95869 274651 95897
rect 274437 95807 274465 95835
rect 274499 95807 274527 95835
rect 274561 95807 274589 95835
rect 274623 95807 274651 95835
rect 274437 95745 274465 95773
rect 274499 95745 274527 95773
rect 274561 95745 274589 95773
rect 274623 95745 274651 95773
rect 274437 86931 274465 86959
rect 274499 86931 274527 86959
rect 274561 86931 274589 86959
rect 274623 86931 274651 86959
rect 274437 86869 274465 86897
rect 274499 86869 274527 86897
rect 274561 86869 274589 86897
rect 274623 86869 274651 86897
rect 274437 86807 274465 86835
rect 274499 86807 274527 86835
rect 274561 86807 274589 86835
rect 274623 86807 274651 86835
rect 274437 86745 274465 86773
rect 274499 86745 274527 86773
rect 274561 86745 274589 86773
rect 274623 86745 274651 86773
rect 274437 77931 274465 77959
rect 274499 77931 274527 77959
rect 274561 77931 274589 77959
rect 274623 77931 274651 77959
rect 274437 77869 274465 77897
rect 274499 77869 274527 77897
rect 274561 77869 274589 77897
rect 274623 77869 274651 77897
rect 274437 77807 274465 77835
rect 274499 77807 274527 77835
rect 274561 77807 274589 77835
rect 274623 77807 274651 77835
rect 274437 77745 274465 77773
rect 274499 77745 274527 77773
rect 274561 77745 274589 77773
rect 274623 77745 274651 77773
rect 274437 68931 274465 68959
rect 274499 68931 274527 68959
rect 274561 68931 274589 68959
rect 274623 68931 274651 68959
rect 274437 68869 274465 68897
rect 274499 68869 274527 68897
rect 274561 68869 274589 68897
rect 274623 68869 274651 68897
rect 274437 68807 274465 68835
rect 274499 68807 274527 68835
rect 274561 68807 274589 68835
rect 274623 68807 274651 68835
rect 274437 68745 274465 68773
rect 274499 68745 274527 68773
rect 274561 68745 274589 68773
rect 274623 68745 274651 68773
rect 274437 59931 274465 59959
rect 274499 59931 274527 59959
rect 274561 59931 274589 59959
rect 274623 59931 274651 59959
rect 274437 59869 274465 59897
rect 274499 59869 274527 59897
rect 274561 59869 274589 59897
rect 274623 59869 274651 59897
rect 274437 59807 274465 59835
rect 274499 59807 274527 59835
rect 274561 59807 274589 59835
rect 274623 59807 274651 59835
rect 274437 59745 274465 59773
rect 274499 59745 274527 59773
rect 274561 59745 274589 59773
rect 274623 59745 274651 59773
rect 274437 50931 274465 50959
rect 274499 50931 274527 50959
rect 274561 50931 274589 50959
rect 274623 50931 274651 50959
rect 274437 50869 274465 50897
rect 274499 50869 274527 50897
rect 274561 50869 274589 50897
rect 274623 50869 274651 50897
rect 274437 50807 274465 50835
rect 274499 50807 274527 50835
rect 274561 50807 274589 50835
rect 274623 50807 274651 50835
rect 274437 50745 274465 50773
rect 274499 50745 274527 50773
rect 274561 50745 274589 50773
rect 274623 50745 274651 50773
rect 274437 41931 274465 41959
rect 274499 41931 274527 41959
rect 274561 41931 274589 41959
rect 274623 41931 274651 41959
rect 274437 41869 274465 41897
rect 274499 41869 274527 41897
rect 274561 41869 274589 41897
rect 274623 41869 274651 41897
rect 274437 41807 274465 41835
rect 274499 41807 274527 41835
rect 274561 41807 274589 41835
rect 274623 41807 274651 41835
rect 274437 41745 274465 41773
rect 274499 41745 274527 41773
rect 274561 41745 274589 41773
rect 274623 41745 274651 41773
rect 274437 32931 274465 32959
rect 274499 32931 274527 32959
rect 274561 32931 274589 32959
rect 274623 32931 274651 32959
rect 274437 32869 274465 32897
rect 274499 32869 274527 32897
rect 274561 32869 274589 32897
rect 274623 32869 274651 32897
rect 274437 32807 274465 32835
rect 274499 32807 274527 32835
rect 274561 32807 274589 32835
rect 274623 32807 274651 32835
rect 274437 32745 274465 32773
rect 274499 32745 274527 32773
rect 274561 32745 274589 32773
rect 274623 32745 274651 32773
rect 274437 23931 274465 23959
rect 274499 23931 274527 23959
rect 274561 23931 274589 23959
rect 274623 23931 274651 23959
rect 274437 23869 274465 23897
rect 274499 23869 274527 23897
rect 274561 23869 274589 23897
rect 274623 23869 274651 23897
rect 274437 23807 274465 23835
rect 274499 23807 274527 23835
rect 274561 23807 274589 23835
rect 274623 23807 274651 23835
rect 274437 23745 274465 23773
rect 274499 23745 274527 23773
rect 274561 23745 274589 23773
rect 274623 23745 274651 23773
rect 274437 14931 274465 14959
rect 274499 14931 274527 14959
rect 274561 14931 274589 14959
rect 274623 14931 274651 14959
rect 274437 14869 274465 14897
rect 274499 14869 274527 14897
rect 274561 14869 274589 14897
rect 274623 14869 274651 14897
rect 274437 14807 274465 14835
rect 274499 14807 274527 14835
rect 274561 14807 274589 14835
rect 274623 14807 274651 14835
rect 274437 14745 274465 14773
rect 274499 14745 274527 14773
rect 274561 14745 274589 14773
rect 274623 14745 274651 14773
rect 274437 5931 274465 5959
rect 274499 5931 274527 5959
rect 274561 5931 274589 5959
rect 274623 5931 274651 5959
rect 274437 5869 274465 5897
rect 274499 5869 274527 5897
rect 274561 5869 274589 5897
rect 274623 5869 274651 5897
rect 274437 5807 274465 5835
rect 274499 5807 274527 5835
rect 274561 5807 274589 5835
rect 274623 5807 274651 5835
rect 274437 5745 274465 5773
rect 274499 5745 274527 5773
rect 274561 5745 274589 5773
rect 274623 5745 274651 5773
rect 274437 396 274465 424
rect 274499 396 274527 424
rect 274561 396 274589 424
rect 274623 396 274651 424
rect 274437 334 274465 362
rect 274499 334 274527 362
rect 274561 334 274589 362
rect 274623 334 274651 362
rect 274437 272 274465 300
rect 274499 272 274527 300
rect 274561 272 274589 300
rect 274623 272 274651 300
rect 274437 210 274465 238
rect 274499 210 274527 238
rect 274561 210 274589 238
rect 274623 210 274651 238
rect 281577 299162 281605 299190
rect 281639 299162 281667 299190
rect 281701 299162 281729 299190
rect 281763 299162 281791 299190
rect 281577 299100 281605 299128
rect 281639 299100 281667 299128
rect 281701 299100 281729 299128
rect 281763 299100 281791 299128
rect 281577 299038 281605 299066
rect 281639 299038 281667 299066
rect 281701 299038 281729 299066
rect 281763 299038 281791 299066
rect 281577 298976 281605 299004
rect 281639 298976 281667 299004
rect 281701 298976 281729 299004
rect 281763 298976 281791 299004
rect 281577 290931 281605 290959
rect 281639 290931 281667 290959
rect 281701 290931 281729 290959
rect 281763 290931 281791 290959
rect 281577 290869 281605 290897
rect 281639 290869 281667 290897
rect 281701 290869 281729 290897
rect 281763 290869 281791 290897
rect 281577 290807 281605 290835
rect 281639 290807 281667 290835
rect 281701 290807 281729 290835
rect 281763 290807 281791 290835
rect 281577 290745 281605 290773
rect 281639 290745 281667 290773
rect 281701 290745 281729 290773
rect 281763 290745 281791 290773
rect 281577 281931 281605 281959
rect 281639 281931 281667 281959
rect 281701 281931 281729 281959
rect 281763 281931 281791 281959
rect 281577 281869 281605 281897
rect 281639 281869 281667 281897
rect 281701 281869 281729 281897
rect 281763 281869 281791 281897
rect 281577 281807 281605 281835
rect 281639 281807 281667 281835
rect 281701 281807 281729 281835
rect 281763 281807 281791 281835
rect 281577 281745 281605 281773
rect 281639 281745 281667 281773
rect 281701 281745 281729 281773
rect 281763 281745 281791 281773
rect 281577 272931 281605 272959
rect 281639 272931 281667 272959
rect 281701 272931 281729 272959
rect 281763 272931 281791 272959
rect 281577 272869 281605 272897
rect 281639 272869 281667 272897
rect 281701 272869 281729 272897
rect 281763 272869 281791 272897
rect 281577 272807 281605 272835
rect 281639 272807 281667 272835
rect 281701 272807 281729 272835
rect 281763 272807 281791 272835
rect 281577 272745 281605 272773
rect 281639 272745 281667 272773
rect 281701 272745 281729 272773
rect 281763 272745 281791 272773
rect 281577 263931 281605 263959
rect 281639 263931 281667 263959
rect 281701 263931 281729 263959
rect 281763 263931 281791 263959
rect 281577 263869 281605 263897
rect 281639 263869 281667 263897
rect 281701 263869 281729 263897
rect 281763 263869 281791 263897
rect 281577 263807 281605 263835
rect 281639 263807 281667 263835
rect 281701 263807 281729 263835
rect 281763 263807 281791 263835
rect 281577 263745 281605 263773
rect 281639 263745 281667 263773
rect 281701 263745 281729 263773
rect 281763 263745 281791 263773
rect 281577 254931 281605 254959
rect 281639 254931 281667 254959
rect 281701 254931 281729 254959
rect 281763 254931 281791 254959
rect 281577 254869 281605 254897
rect 281639 254869 281667 254897
rect 281701 254869 281729 254897
rect 281763 254869 281791 254897
rect 281577 254807 281605 254835
rect 281639 254807 281667 254835
rect 281701 254807 281729 254835
rect 281763 254807 281791 254835
rect 281577 254745 281605 254773
rect 281639 254745 281667 254773
rect 281701 254745 281729 254773
rect 281763 254745 281791 254773
rect 281577 245931 281605 245959
rect 281639 245931 281667 245959
rect 281701 245931 281729 245959
rect 281763 245931 281791 245959
rect 281577 245869 281605 245897
rect 281639 245869 281667 245897
rect 281701 245869 281729 245897
rect 281763 245869 281791 245897
rect 281577 245807 281605 245835
rect 281639 245807 281667 245835
rect 281701 245807 281729 245835
rect 281763 245807 281791 245835
rect 281577 245745 281605 245773
rect 281639 245745 281667 245773
rect 281701 245745 281729 245773
rect 281763 245745 281791 245773
rect 281577 236931 281605 236959
rect 281639 236931 281667 236959
rect 281701 236931 281729 236959
rect 281763 236931 281791 236959
rect 281577 236869 281605 236897
rect 281639 236869 281667 236897
rect 281701 236869 281729 236897
rect 281763 236869 281791 236897
rect 281577 236807 281605 236835
rect 281639 236807 281667 236835
rect 281701 236807 281729 236835
rect 281763 236807 281791 236835
rect 281577 236745 281605 236773
rect 281639 236745 281667 236773
rect 281701 236745 281729 236773
rect 281763 236745 281791 236773
rect 281577 227931 281605 227959
rect 281639 227931 281667 227959
rect 281701 227931 281729 227959
rect 281763 227931 281791 227959
rect 281577 227869 281605 227897
rect 281639 227869 281667 227897
rect 281701 227869 281729 227897
rect 281763 227869 281791 227897
rect 281577 227807 281605 227835
rect 281639 227807 281667 227835
rect 281701 227807 281729 227835
rect 281763 227807 281791 227835
rect 281577 227745 281605 227773
rect 281639 227745 281667 227773
rect 281701 227745 281729 227773
rect 281763 227745 281791 227773
rect 281577 218931 281605 218959
rect 281639 218931 281667 218959
rect 281701 218931 281729 218959
rect 281763 218931 281791 218959
rect 281577 218869 281605 218897
rect 281639 218869 281667 218897
rect 281701 218869 281729 218897
rect 281763 218869 281791 218897
rect 281577 218807 281605 218835
rect 281639 218807 281667 218835
rect 281701 218807 281729 218835
rect 281763 218807 281791 218835
rect 281577 218745 281605 218773
rect 281639 218745 281667 218773
rect 281701 218745 281729 218773
rect 281763 218745 281791 218773
rect 281577 209931 281605 209959
rect 281639 209931 281667 209959
rect 281701 209931 281729 209959
rect 281763 209931 281791 209959
rect 281577 209869 281605 209897
rect 281639 209869 281667 209897
rect 281701 209869 281729 209897
rect 281763 209869 281791 209897
rect 281577 209807 281605 209835
rect 281639 209807 281667 209835
rect 281701 209807 281729 209835
rect 281763 209807 281791 209835
rect 281577 209745 281605 209773
rect 281639 209745 281667 209773
rect 281701 209745 281729 209773
rect 281763 209745 281791 209773
rect 281577 200931 281605 200959
rect 281639 200931 281667 200959
rect 281701 200931 281729 200959
rect 281763 200931 281791 200959
rect 281577 200869 281605 200897
rect 281639 200869 281667 200897
rect 281701 200869 281729 200897
rect 281763 200869 281791 200897
rect 281577 200807 281605 200835
rect 281639 200807 281667 200835
rect 281701 200807 281729 200835
rect 281763 200807 281791 200835
rect 281577 200745 281605 200773
rect 281639 200745 281667 200773
rect 281701 200745 281729 200773
rect 281763 200745 281791 200773
rect 281577 191931 281605 191959
rect 281639 191931 281667 191959
rect 281701 191931 281729 191959
rect 281763 191931 281791 191959
rect 281577 191869 281605 191897
rect 281639 191869 281667 191897
rect 281701 191869 281729 191897
rect 281763 191869 281791 191897
rect 281577 191807 281605 191835
rect 281639 191807 281667 191835
rect 281701 191807 281729 191835
rect 281763 191807 281791 191835
rect 281577 191745 281605 191773
rect 281639 191745 281667 191773
rect 281701 191745 281729 191773
rect 281763 191745 281791 191773
rect 281577 182931 281605 182959
rect 281639 182931 281667 182959
rect 281701 182931 281729 182959
rect 281763 182931 281791 182959
rect 281577 182869 281605 182897
rect 281639 182869 281667 182897
rect 281701 182869 281729 182897
rect 281763 182869 281791 182897
rect 281577 182807 281605 182835
rect 281639 182807 281667 182835
rect 281701 182807 281729 182835
rect 281763 182807 281791 182835
rect 281577 182745 281605 182773
rect 281639 182745 281667 182773
rect 281701 182745 281729 182773
rect 281763 182745 281791 182773
rect 281577 173931 281605 173959
rect 281639 173931 281667 173959
rect 281701 173931 281729 173959
rect 281763 173931 281791 173959
rect 281577 173869 281605 173897
rect 281639 173869 281667 173897
rect 281701 173869 281729 173897
rect 281763 173869 281791 173897
rect 281577 173807 281605 173835
rect 281639 173807 281667 173835
rect 281701 173807 281729 173835
rect 281763 173807 281791 173835
rect 281577 173745 281605 173773
rect 281639 173745 281667 173773
rect 281701 173745 281729 173773
rect 281763 173745 281791 173773
rect 281577 164931 281605 164959
rect 281639 164931 281667 164959
rect 281701 164931 281729 164959
rect 281763 164931 281791 164959
rect 281577 164869 281605 164897
rect 281639 164869 281667 164897
rect 281701 164869 281729 164897
rect 281763 164869 281791 164897
rect 281577 164807 281605 164835
rect 281639 164807 281667 164835
rect 281701 164807 281729 164835
rect 281763 164807 281791 164835
rect 281577 164745 281605 164773
rect 281639 164745 281667 164773
rect 281701 164745 281729 164773
rect 281763 164745 281791 164773
rect 281577 155931 281605 155959
rect 281639 155931 281667 155959
rect 281701 155931 281729 155959
rect 281763 155931 281791 155959
rect 281577 155869 281605 155897
rect 281639 155869 281667 155897
rect 281701 155869 281729 155897
rect 281763 155869 281791 155897
rect 281577 155807 281605 155835
rect 281639 155807 281667 155835
rect 281701 155807 281729 155835
rect 281763 155807 281791 155835
rect 281577 155745 281605 155773
rect 281639 155745 281667 155773
rect 281701 155745 281729 155773
rect 281763 155745 281791 155773
rect 281577 146931 281605 146959
rect 281639 146931 281667 146959
rect 281701 146931 281729 146959
rect 281763 146931 281791 146959
rect 281577 146869 281605 146897
rect 281639 146869 281667 146897
rect 281701 146869 281729 146897
rect 281763 146869 281791 146897
rect 281577 146807 281605 146835
rect 281639 146807 281667 146835
rect 281701 146807 281729 146835
rect 281763 146807 281791 146835
rect 281577 146745 281605 146773
rect 281639 146745 281667 146773
rect 281701 146745 281729 146773
rect 281763 146745 281791 146773
rect 281577 137931 281605 137959
rect 281639 137931 281667 137959
rect 281701 137931 281729 137959
rect 281763 137931 281791 137959
rect 281577 137869 281605 137897
rect 281639 137869 281667 137897
rect 281701 137869 281729 137897
rect 281763 137869 281791 137897
rect 281577 137807 281605 137835
rect 281639 137807 281667 137835
rect 281701 137807 281729 137835
rect 281763 137807 281791 137835
rect 281577 137745 281605 137773
rect 281639 137745 281667 137773
rect 281701 137745 281729 137773
rect 281763 137745 281791 137773
rect 281577 128931 281605 128959
rect 281639 128931 281667 128959
rect 281701 128931 281729 128959
rect 281763 128931 281791 128959
rect 281577 128869 281605 128897
rect 281639 128869 281667 128897
rect 281701 128869 281729 128897
rect 281763 128869 281791 128897
rect 281577 128807 281605 128835
rect 281639 128807 281667 128835
rect 281701 128807 281729 128835
rect 281763 128807 281791 128835
rect 281577 128745 281605 128773
rect 281639 128745 281667 128773
rect 281701 128745 281729 128773
rect 281763 128745 281791 128773
rect 281577 119931 281605 119959
rect 281639 119931 281667 119959
rect 281701 119931 281729 119959
rect 281763 119931 281791 119959
rect 281577 119869 281605 119897
rect 281639 119869 281667 119897
rect 281701 119869 281729 119897
rect 281763 119869 281791 119897
rect 281577 119807 281605 119835
rect 281639 119807 281667 119835
rect 281701 119807 281729 119835
rect 281763 119807 281791 119835
rect 281577 119745 281605 119773
rect 281639 119745 281667 119773
rect 281701 119745 281729 119773
rect 281763 119745 281791 119773
rect 281577 110931 281605 110959
rect 281639 110931 281667 110959
rect 281701 110931 281729 110959
rect 281763 110931 281791 110959
rect 281577 110869 281605 110897
rect 281639 110869 281667 110897
rect 281701 110869 281729 110897
rect 281763 110869 281791 110897
rect 281577 110807 281605 110835
rect 281639 110807 281667 110835
rect 281701 110807 281729 110835
rect 281763 110807 281791 110835
rect 281577 110745 281605 110773
rect 281639 110745 281667 110773
rect 281701 110745 281729 110773
rect 281763 110745 281791 110773
rect 281577 101931 281605 101959
rect 281639 101931 281667 101959
rect 281701 101931 281729 101959
rect 281763 101931 281791 101959
rect 281577 101869 281605 101897
rect 281639 101869 281667 101897
rect 281701 101869 281729 101897
rect 281763 101869 281791 101897
rect 281577 101807 281605 101835
rect 281639 101807 281667 101835
rect 281701 101807 281729 101835
rect 281763 101807 281791 101835
rect 281577 101745 281605 101773
rect 281639 101745 281667 101773
rect 281701 101745 281729 101773
rect 281763 101745 281791 101773
rect 281577 92931 281605 92959
rect 281639 92931 281667 92959
rect 281701 92931 281729 92959
rect 281763 92931 281791 92959
rect 281577 92869 281605 92897
rect 281639 92869 281667 92897
rect 281701 92869 281729 92897
rect 281763 92869 281791 92897
rect 281577 92807 281605 92835
rect 281639 92807 281667 92835
rect 281701 92807 281729 92835
rect 281763 92807 281791 92835
rect 281577 92745 281605 92773
rect 281639 92745 281667 92773
rect 281701 92745 281729 92773
rect 281763 92745 281791 92773
rect 281577 83931 281605 83959
rect 281639 83931 281667 83959
rect 281701 83931 281729 83959
rect 281763 83931 281791 83959
rect 281577 83869 281605 83897
rect 281639 83869 281667 83897
rect 281701 83869 281729 83897
rect 281763 83869 281791 83897
rect 281577 83807 281605 83835
rect 281639 83807 281667 83835
rect 281701 83807 281729 83835
rect 281763 83807 281791 83835
rect 281577 83745 281605 83773
rect 281639 83745 281667 83773
rect 281701 83745 281729 83773
rect 281763 83745 281791 83773
rect 281577 74931 281605 74959
rect 281639 74931 281667 74959
rect 281701 74931 281729 74959
rect 281763 74931 281791 74959
rect 281577 74869 281605 74897
rect 281639 74869 281667 74897
rect 281701 74869 281729 74897
rect 281763 74869 281791 74897
rect 281577 74807 281605 74835
rect 281639 74807 281667 74835
rect 281701 74807 281729 74835
rect 281763 74807 281791 74835
rect 281577 74745 281605 74773
rect 281639 74745 281667 74773
rect 281701 74745 281729 74773
rect 281763 74745 281791 74773
rect 281577 65931 281605 65959
rect 281639 65931 281667 65959
rect 281701 65931 281729 65959
rect 281763 65931 281791 65959
rect 281577 65869 281605 65897
rect 281639 65869 281667 65897
rect 281701 65869 281729 65897
rect 281763 65869 281791 65897
rect 281577 65807 281605 65835
rect 281639 65807 281667 65835
rect 281701 65807 281729 65835
rect 281763 65807 281791 65835
rect 281577 65745 281605 65773
rect 281639 65745 281667 65773
rect 281701 65745 281729 65773
rect 281763 65745 281791 65773
rect 281577 56931 281605 56959
rect 281639 56931 281667 56959
rect 281701 56931 281729 56959
rect 281763 56931 281791 56959
rect 281577 56869 281605 56897
rect 281639 56869 281667 56897
rect 281701 56869 281729 56897
rect 281763 56869 281791 56897
rect 281577 56807 281605 56835
rect 281639 56807 281667 56835
rect 281701 56807 281729 56835
rect 281763 56807 281791 56835
rect 281577 56745 281605 56773
rect 281639 56745 281667 56773
rect 281701 56745 281729 56773
rect 281763 56745 281791 56773
rect 281577 47931 281605 47959
rect 281639 47931 281667 47959
rect 281701 47931 281729 47959
rect 281763 47931 281791 47959
rect 281577 47869 281605 47897
rect 281639 47869 281667 47897
rect 281701 47869 281729 47897
rect 281763 47869 281791 47897
rect 281577 47807 281605 47835
rect 281639 47807 281667 47835
rect 281701 47807 281729 47835
rect 281763 47807 281791 47835
rect 281577 47745 281605 47773
rect 281639 47745 281667 47773
rect 281701 47745 281729 47773
rect 281763 47745 281791 47773
rect 281577 38931 281605 38959
rect 281639 38931 281667 38959
rect 281701 38931 281729 38959
rect 281763 38931 281791 38959
rect 281577 38869 281605 38897
rect 281639 38869 281667 38897
rect 281701 38869 281729 38897
rect 281763 38869 281791 38897
rect 281577 38807 281605 38835
rect 281639 38807 281667 38835
rect 281701 38807 281729 38835
rect 281763 38807 281791 38835
rect 281577 38745 281605 38773
rect 281639 38745 281667 38773
rect 281701 38745 281729 38773
rect 281763 38745 281791 38773
rect 281577 29931 281605 29959
rect 281639 29931 281667 29959
rect 281701 29931 281729 29959
rect 281763 29931 281791 29959
rect 281577 29869 281605 29897
rect 281639 29869 281667 29897
rect 281701 29869 281729 29897
rect 281763 29869 281791 29897
rect 281577 29807 281605 29835
rect 281639 29807 281667 29835
rect 281701 29807 281729 29835
rect 281763 29807 281791 29835
rect 281577 29745 281605 29773
rect 281639 29745 281667 29773
rect 281701 29745 281729 29773
rect 281763 29745 281791 29773
rect 281577 20931 281605 20959
rect 281639 20931 281667 20959
rect 281701 20931 281729 20959
rect 281763 20931 281791 20959
rect 281577 20869 281605 20897
rect 281639 20869 281667 20897
rect 281701 20869 281729 20897
rect 281763 20869 281791 20897
rect 281577 20807 281605 20835
rect 281639 20807 281667 20835
rect 281701 20807 281729 20835
rect 281763 20807 281791 20835
rect 281577 20745 281605 20773
rect 281639 20745 281667 20773
rect 281701 20745 281729 20773
rect 281763 20745 281791 20773
rect 281577 11931 281605 11959
rect 281639 11931 281667 11959
rect 281701 11931 281729 11959
rect 281763 11931 281791 11959
rect 281577 11869 281605 11897
rect 281639 11869 281667 11897
rect 281701 11869 281729 11897
rect 281763 11869 281791 11897
rect 281577 11807 281605 11835
rect 281639 11807 281667 11835
rect 281701 11807 281729 11835
rect 281763 11807 281791 11835
rect 281577 11745 281605 11773
rect 281639 11745 281667 11773
rect 281701 11745 281729 11773
rect 281763 11745 281791 11773
rect 281577 2931 281605 2959
rect 281639 2931 281667 2959
rect 281701 2931 281729 2959
rect 281763 2931 281791 2959
rect 281577 2869 281605 2897
rect 281639 2869 281667 2897
rect 281701 2869 281729 2897
rect 281763 2869 281791 2897
rect 281577 2807 281605 2835
rect 281639 2807 281667 2835
rect 281701 2807 281729 2835
rect 281763 2807 281791 2835
rect 281577 2745 281605 2773
rect 281639 2745 281667 2773
rect 281701 2745 281729 2773
rect 281763 2745 281791 2773
rect 281577 876 281605 904
rect 281639 876 281667 904
rect 281701 876 281729 904
rect 281763 876 281791 904
rect 281577 814 281605 842
rect 281639 814 281667 842
rect 281701 814 281729 842
rect 281763 814 281791 842
rect 281577 752 281605 780
rect 281639 752 281667 780
rect 281701 752 281729 780
rect 281763 752 281791 780
rect 281577 690 281605 718
rect 281639 690 281667 718
rect 281701 690 281729 718
rect 281763 690 281791 718
rect 283437 299642 283465 299670
rect 283499 299642 283527 299670
rect 283561 299642 283589 299670
rect 283623 299642 283651 299670
rect 283437 299580 283465 299608
rect 283499 299580 283527 299608
rect 283561 299580 283589 299608
rect 283623 299580 283651 299608
rect 283437 299518 283465 299546
rect 283499 299518 283527 299546
rect 283561 299518 283589 299546
rect 283623 299518 283651 299546
rect 283437 299456 283465 299484
rect 283499 299456 283527 299484
rect 283561 299456 283589 299484
rect 283623 299456 283651 299484
rect 283437 293931 283465 293959
rect 283499 293931 283527 293959
rect 283561 293931 283589 293959
rect 283623 293931 283651 293959
rect 283437 293869 283465 293897
rect 283499 293869 283527 293897
rect 283561 293869 283589 293897
rect 283623 293869 283651 293897
rect 283437 293807 283465 293835
rect 283499 293807 283527 293835
rect 283561 293807 283589 293835
rect 283623 293807 283651 293835
rect 283437 293745 283465 293773
rect 283499 293745 283527 293773
rect 283561 293745 283589 293773
rect 283623 293745 283651 293773
rect 283437 284931 283465 284959
rect 283499 284931 283527 284959
rect 283561 284931 283589 284959
rect 283623 284931 283651 284959
rect 283437 284869 283465 284897
rect 283499 284869 283527 284897
rect 283561 284869 283589 284897
rect 283623 284869 283651 284897
rect 283437 284807 283465 284835
rect 283499 284807 283527 284835
rect 283561 284807 283589 284835
rect 283623 284807 283651 284835
rect 283437 284745 283465 284773
rect 283499 284745 283527 284773
rect 283561 284745 283589 284773
rect 283623 284745 283651 284773
rect 283437 275931 283465 275959
rect 283499 275931 283527 275959
rect 283561 275931 283589 275959
rect 283623 275931 283651 275959
rect 283437 275869 283465 275897
rect 283499 275869 283527 275897
rect 283561 275869 283589 275897
rect 283623 275869 283651 275897
rect 283437 275807 283465 275835
rect 283499 275807 283527 275835
rect 283561 275807 283589 275835
rect 283623 275807 283651 275835
rect 283437 275745 283465 275773
rect 283499 275745 283527 275773
rect 283561 275745 283589 275773
rect 283623 275745 283651 275773
rect 283437 266931 283465 266959
rect 283499 266931 283527 266959
rect 283561 266931 283589 266959
rect 283623 266931 283651 266959
rect 283437 266869 283465 266897
rect 283499 266869 283527 266897
rect 283561 266869 283589 266897
rect 283623 266869 283651 266897
rect 283437 266807 283465 266835
rect 283499 266807 283527 266835
rect 283561 266807 283589 266835
rect 283623 266807 283651 266835
rect 283437 266745 283465 266773
rect 283499 266745 283527 266773
rect 283561 266745 283589 266773
rect 283623 266745 283651 266773
rect 283437 257931 283465 257959
rect 283499 257931 283527 257959
rect 283561 257931 283589 257959
rect 283623 257931 283651 257959
rect 283437 257869 283465 257897
rect 283499 257869 283527 257897
rect 283561 257869 283589 257897
rect 283623 257869 283651 257897
rect 283437 257807 283465 257835
rect 283499 257807 283527 257835
rect 283561 257807 283589 257835
rect 283623 257807 283651 257835
rect 283437 257745 283465 257773
rect 283499 257745 283527 257773
rect 283561 257745 283589 257773
rect 283623 257745 283651 257773
rect 283437 248931 283465 248959
rect 283499 248931 283527 248959
rect 283561 248931 283589 248959
rect 283623 248931 283651 248959
rect 283437 248869 283465 248897
rect 283499 248869 283527 248897
rect 283561 248869 283589 248897
rect 283623 248869 283651 248897
rect 283437 248807 283465 248835
rect 283499 248807 283527 248835
rect 283561 248807 283589 248835
rect 283623 248807 283651 248835
rect 283437 248745 283465 248773
rect 283499 248745 283527 248773
rect 283561 248745 283589 248773
rect 283623 248745 283651 248773
rect 283437 239931 283465 239959
rect 283499 239931 283527 239959
rect 283561 239931 283589 239959
rect 283623 239931 283651 239959
rect 283437 239869 283465 239897
rect 283499 239869 283527 239897
rect 283561 239869 283589 239897
rect 283623 239869 283651 239897
rect 283437 239807 283465 239835
rect 283499 239807 283527 239835
rect 283561 239807 283589 239835
rect 283623 239807 283651 239835
rect 283437 239745 283465 239773
rect 283499 239745 283527 239773
rect 283561 239745 283589 239773
rect 283623 239745 283651 239773
rect 283437 230931 283465 230959
rect 283499 230931 283527 230959
rect 283561 230931 283589 230959
rect 283623 230931 283651 230959
rect 283437 230869 283465 230897
rect 283499 230869 283527 230897
rect 283561 230869 283589 230897
rect 283623 230869 283651 230897
rect 283437 230807 283465 230835
rect 283499 230807 283527 230835
rect 283561 230807 283589 230835
rect 283623 230807 283651 230835
rect 283437 230745 283465 230773
rect 283499 230745 283527 230773
rect 283561 230745 283589 230773
rect 283623 230745 283651 230773
rect 283437 221931 283465 221959
rect 283499 221931 283527 221959
rect 283561 221931 283589 221959
rect 283623 221931 283651 221959
rect 283437 221869 283465 221897
rect 283499 221869 283527 221897
rect 283561 221869 283589 221897
rect 283623 221869 283651 221897
rect 283437 221807 283465 221835
rect 283499 221807 283527 221835
rect 283561 221807 283589 221835
rect 283623 221807 283651 221835
rect 283437 221745 283465 221773
rect 283499 221745 283527 221773
rect 283561 221745 283589 221773
rect 283623 221745 283651 221773
rect 283437 212931 283465 212959
rect 283499 212931 283527 212959
rect 283561 212931 283589 212959
rect 283623 212931 283651 212959
rect 283437 212869 283465 212897
rect 283499 212869 283527 212897
rect 283561 212869 283589 212897
rect 283623 212869 283651 212897
rect 283437 212807 283465 212835
rect 283499 212807 283527 212835
rect 283561 212807 283589 212835
rect 283623 212807 283651 212835
rect 283437 212745 283465 212773
rect 283499 212745 283527 212773
rect 283561 212745 283589 212773
rect 283623 212745 283651 212773
rect 283437 203931 283465 203959
rect 283499 203931 283527 203959
rect 283561 203931 283589 203959
rect 283623 203931 283651 203959
rect 283437 203869 283465 203897
rect 283499 203869 283527 203897
rect 283561 203869 283589 203897
rect 283623 203869 283651 203897
rect 283437 203807 283465 203835
rect 283499 203807 283527 203835
rect 283561 203807 283589 203835
rect 283623 203807 283651 203835
rect 283437 203745 283465 203773
rect 283499 203745 283527 203773
rect 283561 203745 283589 203773
rect 283623 203745 283651 203773
rect 283437 194931 283465 194959
rect 283499 194931 283527 194959
rect 283561 194931 283589 194959
rect 283623 194931 283651 194959
rect 283437 194869 283465 194897
rect 283499 194869 283527 194897
rect 283561 194869 283589 194897
rect 283623 194869 283651 194897
rect 283437 194807 283465 194835
rect 283499 194807 283527 194835
rect 283561 194807 283589 194835
rect 283623 194807 283651 194835
rect 283437 194745 283465 194773
rect 283499 194745 283527 194773
rect 283561 194745 283589 194773
rect 283623 194745 283651 194773
rect 283437 185931 283465 185959
rect 283499 185931 283527 185959
rect 283561 185931 283589 185959
rect 283623 185931 283651 185959
rect 283437 185869 283465 185897
rect 283499 185869 283527 185897
rect 283561 185869 283589 185897
rect 283623 185869 283651 185897
rect 283437 185807 283465 185835
rect 283499 185807 283527 185835
rect 283561 185807 283589 185835
rect 283623 185807 283651 185835
rect 283437 185745 283465 185773
rect 283499 185745 283527 185773
rect 283561 185745 283589 185773
rect 283623 185745 283651 185773
rect 283437 176931 283465 176959
rect 283499 176931 283527 176959
rect 283561 176931 283589 176959
rect 283623 176931 283651 176959
rect 283437 176869 283465 176897
rect 283499 176869 283527 176897
rect 283561 176869 283589 176897
rect 283623 176869 283651 176897
rect 283437 176807 283465 176835
rect 283499 176807 283527 176835
rect 283561 176807 283589 176835
rect 283623 176807 283651 176835
rect 283437 176745 283465 176773
rect 283499 176745 283527 176773
rect 283561 176745 283589 176773
rect 283623 176745 283651 176773
rect 283437 167931 283465 167959
rect 283499 167931 283527 167959
rect 283561 167931 283589 167959
rect 283623 167931 283651 167959
rect 283437 167869 283465 167897
rect 283499 167869 283527 167897
rect 283561 167869 283589 167897
rect 283623 167869 283651 167897
rect 283437 167807 283465 167835
rect 283499 167807 283527 167835
rect 283561 167807 283589 167835
rect 283623 167807 283651 167835
rect 283437 167745 283465 167773
rect 283499 167745 283527 167773
rect 283561 167745 283589 167773
rect 283623 167745 283651 167773
rect 283437 158931 283465 158959
rect 283499 158931 283527 158959
rect 283561 158931 283589 158959
rect 283623 158931 283651 158959
rect 283437 158869 283465 158897
rect 283499 158869 283527 158897
rect 283561 158869 283589 158897
rect 283623 158869 283651 158897
rect 283437 158807 283465 158835
rect 283499 158807 283527 158835
rect 283561 158807 283589 158835
rect 283623 158807 283651 158835
rect 283437 158745 283465 158773
rect 283499 158745 283527 158773
rect 283561 158745 283589 158773
rect 283623 158745 283651 158773
rect 283437 149931 283465 149959
rect 283499 149931 283527 149959
rect 283561 149931 283589 149959
rect 283623 149931 283651 149959
rect 283437 149869 283465 149897
rect 283499 149869 283527 149897
rect 283561 149869 283589 149897
rect 283623 149869 283651 149897
rect 283437 149807 283465 149835
rect 283499 149807 283527 149835
rect 283561 149807 283589 149835
rect 283623 149807 283651 149835
rect 283437 149745 283465 149773
rect 283499 149745 283527 149773
rect 283561 149745 283589 149773
rect 283623 149745 283651 149773
rect 283437 140931 283465 140959
rect 283499 140931 283527 140959
rect 283561 140931 283589 140959
rect 283623 140931 283651 140959
rect 283437 140869 283465 140897
rect 283499 140869 283527 140897
rect 283561 140869 283589 140897
rect 283623 140869 283651 140897
rect 283437 140807 283465 140835
rect 283499 140807 283527 140835
rect 283561 140807 283589 140835
rect 283623 140807 283651 140835
rect 283437 140745 283465 140773
rect 283499 140745 283527 140773
rect 283561 140745 283589 140773
rect 283623 140745 283651 140773
rect 283437 131931 283465 131959
rect 283499 131931 283527 131959
rect 283561 131931 283589 131959
rect 283623 131931 283651 131959
rect 283437 131869 283465 131897
rect 283499 131869 283527 131897
rect 283561 131869 283589 131897
rect 283623 131869 283651 131897
rect 283437 131807 283465 131835
rect 283499 131807 283527 131835
rect 283561 131807 283589 131835
rect 283623 131807 283651 131835
rect 283437 131745 283465 131773
rect 283499 131745 283527 131773
rect 283561 131745 283589 131773
rect 283623 131745 283651 131773
rect 283437 122931 283465 122959
rect 283499 122931 283527 122959
rect 283561 122931 283589 122959
rect 283623 122931 283651 122959
rect 283437 122869 283465 122897
rect 283499 122869 283527 122897
rect 283561 122869 283589 122897
rect 283623 122869 283651 122897
rect 283437 122807 283465 122835
rect 283499 122807 283527 122835
rect 283561 122807 283589 122835
rect 283623 122807 283651 122835
rect 283437 122745 283465 122773
rect 283499 122745 283527 122773
rect 283561 122745 283589 122773
rect 283623 122745 283651 122773
rect 283437 113931 283465 113959
rect 283499 113931 283527 113959
rect 283561 113931 283589 113959
rect 283623 113931 283651 113959
rect 283437 113869 283465 113897
rect 283499 113869 283527 113897
rect 283561 113869 283589 113897
rect 283623 113869 283651 113897
rect 283437 113807 283465 113835
rect 283499 113807 283527 113835
rect 283561 113807 283589 113835
rect 283623 113807 283651 113835
rect 283437 113745 283465 113773
rect 283499 113745 283527 113773
rect 283561 113745 283589 113773
rect 283623 113745 283651 113773
rect 283437 104931 283465 104959
rect 283499 104931 283527 104959
rect 283561 104931 283589 104959
rect 283623 104931 283651 104959
rect 283437 104869 283465 104897
rect 283499 104869 283527 104897
rect 283561 104869 283589 104897
rect 283623 104869 283651 104897
rect 283437 104807 283465 104835
rect 283499 104807 283527 104835
rect 283561 104807 283589 104835
rect 283623 104807 283651 104835
rect 283437 104745 283465 104773
rect 283499 104745 283527 104773
rect 283561 104745 283589 104773
rect 283623 104745 283651 104773
rect 283437 95931 283465 95959
rect 283499 95931 283527 95959
rect 283561 95931 283589 95959
rect 283623 95931 283651 95959
rect 283437 95869 283465 95897
rect 283499 95869 283527 95897
rect 283561 95869 283589 95897
rect 283623 95869 283651 95897
rect 283437 95807 283465 95835
rect 283499 95807 283527 95835
rect 283561 95807 283589 95835
rect 283623 95807 283651 95835
rect 283437 95745 283465 95773
rect 283499 95745 283527 95773
rect 283561 95745 283589 95773
rect 283623 95745 283651 95773
rect 283437 86931 283465 86959
rect 283499 86931 283527 86959
rect 283561 86931 283589 86959
rect 283623 86931 283651 86959
rect 283437 86869 283465 86897
rect 283499 86869 283527 86897
rect 283561 86869 283589 86897
rect 283623 86869 283651 86897
rect 283437 86807 283465 86835
rect 283499 86807 283527 86835
rect 283561 86807 283589 86835
rect 283623 86807 283651 86835
rect 283437 86745 283465 86773
rect 283499 86745 283527 86773
rect 283561 86745 283589 86773
rect 283623 86745 283651 86773
rect 283437 77931 283465 77959
rect 283499 77931 283527 77959
rect 283561 77931 283589 77959
rect 283623 77931 283651 77959
rect 283437 77869 283465 77897
rect 283499 77869 283527 77897
rect 283561 77869 283589 77897
rect 283623 77869 283651 77897
rect 283437 77807 283465 77835
rect 283499 77807 283527 77835
rect 283561 77807 283589 77835
rect 283623 77807 283651 77835
rect 283437 77745 283465 77773
rect 283499 77745 283527 77773
rect 283561 77745 283589 77773
rect 283623 77745 283651 77773
rect 283437 68931 283465 68959
rect 283499 68931 283527 68959
rect 283561 68931 283589 68959
rect 283623 68931 283651 68959
rect 283437 68869 283465 68897
rect 283499 68869 283527 68897
rect 283561 68869 283589 68897
rect 283623 68869 283651 68897
rect 283437 68807 283465 68835
rect 283499 68807 283527 68835
rect 283561 68807 283589 68835
rect 283623 68807 283651 68835
rect 283437 68745 283465 68773
rect 283499 68745 283527 68773
rect 283561 68745 283589 68773
rect 283623 68745 283651 68773
rect 283437 59931 283465 59959
rect 283499 59931 283527 59959
rect 283561 59931 283589 59959
rect 283623 59931 283651 59959
rect 283437 59869 283465 59897
rect 283499 59869 283527 59897
rect 283561 59869 283589 59897
rect 283623 59869 283651 59897
rect 283437 59807 283465 59835
rect 283499 59807 283527 59835
rect 283561 59807 283589 59835
rect 283623 59807 283651 59835
rect 283437 59745 283465 59773
rect 283499 59745 283527 59773
rect 283561 59745 283589 59773
rect 283623 59745 283651 59773
rect 283437 50931 283465 50959
rect 283499 50931 283527 50959
rect 283561 50931 283589 50959
rect 283623 50931 283651 50959
rect 283437 50869 283465 50897
rect 283499 50869 283527 50897
rect 283561 50869 283589 50897
rect 283623 50869 283651 50897
rect 283437 50807 283465 50835
rect 283499 50807 283527 50835
rect 283561 50807 283589 50835
rect 283623 50807 283651 50835
rect 283437 50745 283465 50773
rect 283499 50745 283527 50773
rect 283561 50745 283589 50773
rect 283623 50745 283651 50773
rect 283437 41931 283465 41959
rect 283499 41931 283527 41959
rect 283561 41931 283589 41959
rect 283623 41931 283651 41959
rect 283437 41869 283465 41897
rect 283499 41869 283527 41897
rect 283561 41869 283589 41897
rect 283623 41869 283651 41897
rect 283437 41807 283465 41835
rect 283499 41807 283527 41835
rect 283561 41807 283589 41835
rect 283623 41807 283651 41835
rect 283437 41745 283465 41773
rect 283499 41745 283527 41773
rect 283561 41745 283589 41773
rect 283623 41745 283651 41773
rect 283437 32931 283465 32959
rect 283499 32931 283527 32959
rect 283561 32931 283589 32959
rect 283623 32931 283651 32959
rect 283437 32869 283465 32897
rect 283499 32869 283527 32897
rect 283561 32869 283589 32897
rect 283623 32869 283651 32897
rect 283437 32807 283465 32835
rect 283499 32807 283527 32835
rect 283561 32807 283589 32835
rect 283623 32807 283651 32835
rect 283437 32745 283465 32773
rect 283499 32745 283527 32773
rect 283561 32745 283589 32773
rect 283623 32745 283651 32773
rect 283437 23931 283465 23959
rect 283499 23931 283527 23959
rect 283561 23931 283589 23959
rect 283623 23931 283651 23959
rect 283437 23869 283465 23897
rect 283499 23869 283527 23897
rect 283561 23869 283589 23897
rect 283623 23869 283651 23897
rect 283437 23807 283465 23835
rect 283499 23807 283527 23835
rect 283561 23807 283589 23835
rect 283623 23807 283651 23835
rect 283437 23745 283465 23773
rect 283499 23745 283527 23773
rect 283561 23745 283589 23773
rect 283623 23745 283651 23773
rect 283437 14931 283465 14959
rect 283499 14931 283527 14959
rect 283561 14931 283589 14959
rect 283623 14931 283651 14959
rect 283437 14869 283465 14897
rect 283499 14869 283527 14897
rect 283561 14869 283589 14897
rect 283623 14869 283651 14897
rect 283437 14807 283465 14835
rect 283499 14807 283527 14835
rect 283561 14807 283589 14835
rect 283623 14807 283651 14835
rect 283437 14745 283465 14773
rect 283499 14745 283527 14773
rect 283561 14745 283589 14773
rect 283623 14745 283651 14773
rect 283437 5931 283465 5959
rect 283499 5931 283527 5959
rect 283561 5931 283589 5959
rect 283623 5931 283651 5959
rect 283437 5869 283465 5897
rect 283499 5869 283527 5897
rect 283561 5869 283589 5897
rect 283623 5869 283651 5897
rect 283437 5807 283465 5835
rect 283499 5807 283527 5835
rect 283561 5807 283589 5835
rect 283623 5807 283651 5835
rect 283437 5745 283465 5773
rect 283499 5745 283527 5773
rect 283561 5745 283589 5773
rect 283623 5745 283651 5773
rect 283437 396 283465 424
rect 283499 396 283527 424
rect 283561 396 283589 424
rect 283623 396 283651 424
rect 283437 334 283465 362
rect 283499 334 283527 362
rect 283561 334 283589 362
rect 283623 334 283651 362
rect 283437 272 283465 300
rect 283499 272 283527 300
rect 283561 272 283589 300
rect 283623 272 283651 300
rect 283437 210 283465 238
rect 283499 210 283527 238
rect 283561 210 283589 238
rect 283623 210 283651 238
rect 290577 299162 290605 299190
rect 290639 299162 290667 299190
rect 290701 299162 290729 299190
rect 290763 299162 290791 299190
rect 290577 299100 290605 299128
rect 290639 299100 290667 299128
rect 290701 299100 290729 299128
rect 290763 299100 290791 299128
rect 290577 299038 290605 299066
rect 290639 299038 290667 299066
rect 290701 299038 290729 299066
rect 290763 299038 290791 299066
rect 290577 298976 290605 299004
rect 290639 298976 290667 299004
rect 290701 298976 290729 299004
rect 290763 298976 290791 299004
rect 290577 290931 290605 290959
rect 290639 290931 290667 290959
rect 290701 290931 290729 290959
rect 290763 290931 290791 290959
rect 290577 290869 290605 290897
rect 290639 290869 290667 290897
rect 290701 290869 290729 290897
rect 290763 290869 290791 290897
rect 290577 290807 290605 290835
rect 290639 290807 290667 290835
rect 290701 290807 290729 290835
rect 290763 290807 290791 290835
rect 290577 290745 290605 290773
rect 290639 290745 290667 290773
rect 290701 290745 290729 290773
rect 290763 290745 290791 290773
rect 290577 281931 290605 281959
rect 290639 281931 290667 281959
rect 290701 281931 290729 281959
rect 290763 281931 290791 281959
rect 290577 281869 290605 281897
rect 290639 281869 290667 281897
rect 290701 281869 290729 281897
rect 290763 281869 290791 281897
rect 290577 281807 290605 281835
rect 290639 281807 290667 281835
rect 290701 281807 290729 281835
rect 290763 281807 290791 281835
rect 290577 281745 290605 281773
rect 290639 281745 290667 281773
rect 290701 281745 290729 281773
rect 290763 281745 290791 281773
rect 290577 272931 290605 272959
rect 290639 272931 290667 272959
rect 290701 272931 290729 272959
rect 290763 272931 290791 272959
rect 290577 272869 290605 272897
rect 290639 272869 290667 272897
rect 290701 272869 290729 272897
rect 290763 272869 290791 272897
rect 290577 272807 290605 272835
rect 290639 272807 290667 272835
rect 290701 272807 290729 272835
rect 290763 272807 290791 272835
rect 290577 272745 290605 272773
rect 290639 272745 290667 272773
rect 290701 272745 290729 272773
rect 290763 272745 290791 272773
rect 290577 263931 290605 263959
rect 290639 263931 290667 263959
rect 290701 263931 290729 263959
rect 290763 263931 290791 263959
rect 290577 263869 290605 263897
rect 290639 263869 290667 263897
rect 290701 263869 290729 263897
rect 290763 263869 290791 263897
rect 290577 263807 290605 263835
rect 290639 263807 290667 263835
rect 290701 263807 290729 263835
rect 290763 263807 290791 263835
rect 290577 263745 290605 263773
rect 290639 263745 290667 263773
rect 290701 263745 290729 263773
rect 290763 263745 290791 263773
rect 290577 254931 290605 254959
rect 290639 254931 290667 254959
rect 290701 254931 290729 254959
rect 290763 254931 290791 254959
rect 290577 254869 290605 254897
rect 290639 254869 290667 254897
rect 290701 254869 290729 254897
rect 290763 254869 290791 254897
rect 290577 254807 290605 254835
rect 290639 254807 290667 254835
rect 290701 254807 290729 254835
rect 290763 254807 290791 254835
rect 290577 254745 290605 254773
rect 290639 254745 290667 254773
rect 290701 254745 290729 254773
rect 290763 254745 290791 254773
rect 290577 245931 290605 245959
rect 290639 245931 290667 245959
rect 290701 245931 290729 245959
rect 290763 245931 290791 245959
rect 290577 245869 290605 245897
rect 290639 245869 290667 245897
rect 290701 245869 290729 245897
rect 290763 245869 290791 245897
rect 290577 245807 290605 245835
rect 290639 245807 290667 245835
rect 290701 245807 290729 245835
rect 290763 245807 290791 245835
rect 290577 245745 290605 245773
rect 290639 245745 290667 245773
rect 290701 245745 290729 245773
rect 290763 245745 290791 245773
rect 290577 236931 290605 236959
rect 290639 236931 290667 236959
rect 290701 236931 290729 236959
rect 290763 236931 290791 236959
rect 290577 236869 290605 236897
rect 290639 236869 290667 236897
rect 290701 236869 290729 236897
rect 290763 236869 290791 236897
rect 290577 236807 290605 236835
rect 290639 236807 290667 236835
rect 290701 236807 290729 236835
rect 290763 236807 290791 236835
rect 290577 236745 290605 236773
rect 290639 236745 290667 236773
rect 290701 236745 290729 236773
rect 290763 236745 290791 236773
rect 290577 227931 290605 227959
rect 290639 227931 290667 227959
rect 290701 227931 290729 227959
rect 290763 227931 290791 227959
rect 290577 227869 290605 227897
rect 290639 227869 290667 227897
rect 290701 227869 290729 227897
rect 290763 227869 290791 227897
rect 290577 227807 290605 227835
rect 290639 227807 290667 227835
rect 290701 227807 290729 227835
rect 290763 227807 290791 227835
rect 290577 227745 290605 227773
rect 290639 227745 290667 227773
rect 290701 227745 290729 227773
rect 290763 227745 290791 227773
rect 290577 218931 290605 218959
rect 290639 218931 290667 218959
rect 290701 218931 290729 218959
rect 290763 218931 290791 218959
rect 290577 218869 290605 218897
rect 290639 218869 290667 218897
rect 290701 218869 290729 218897
rect 290763 218869 290791 218897
rect 290577 218807 290605 218835
rect 290639 218807 290667 218835
rect 290701 218807 290729 218835
rect 290763 218807 290791 218835
rect 290577 218745 290605 218773
rect 290639 218745 290667 218773
rect 290701 218745 290729 218773
rect 290763 218745 290791 218773
rect 290577 209931 290605 209959
rect 290639 209931 290667 209959
rect 290701 209931 290729 209959
rect 290763 209931 290791 209959
rect 290577 209869 290605 209897
rect 290639 209869 290667 209897
rect 290701 209869 290729 209897
rect 290763 209869 290791 209897
rect 290577 209807 290605 209835
rect 290639 209807 290667 209835
rect 290701 209807 290729 209835
rect 290763 209807 290791 209835
rect 290577 209745 290605 209773
rect 290639 209745 290667 209773
rect 290701 209745 290729 209773
rect 290763 209745 290791 209773
rect 290577 200931 290605 200959
rect 290639 200931 290667 200959
rect 290701 200931 290729 200959
rect 290763 200931 290791 200959
rect 290577 200869 290605 200897
rect 290639 200869 290667 200897
rect 290701 200869 290729 200897
rect 290763 200869 290791 200897
rect 290577 200807 290605 200835
rect 290639 200807 290667 200835
rect 290701 200807 290729 200835
rect 290763 200807 290791 200835
rect 290577 200745 290605 200773
rect 290639 200745 290667 200773
rect 290701 200745 290729 200773
rect 290763 200745 290791 200773
rect 290577 191931 290605 191959
rect 290639 191931 290667 191959
rect 290701 191931 290729 191959
rect 290763 191931 290791 191959
rect 290577 191869 290605 191897
rect 290639 191869 290667 191897
rect 290701 191869 290729 191897
rect 290763 191869 290791 191897
rect 290577 191807 290605 191835
rect 290639 191807 290667 191835
rect 290701 191807 290729 191835
rect 290763 191807 290791 191835
rect 290577 191745 290605 191773
rect 290639 191745 290667 191773
rect 290701 191745 290729 191773
rect 290763 191745 290791 191773
rect 290577 182931 290605 182959
rect 290639 182931 290667 182959
rect 290701 182931 290729 182959
rect 290763 182931 290791 182959
rect 290577 182869 290605 182897
rect 290639 182869 290667 182897
rect 290701 182869 290729 182897
rect 290763 182869 290791 182897
rect 290577 182807 290605 182835
rect 290639 182807 290667 182835
rect 290701 182807 290729 182835
rect 290763 182807 290791 182835
rect 290577 182745 290605 182773
rect 290639 182745 290667 182773
rect 290701 182745 290729 182773
rect 290763 182745 290791 182773
rect 290577 173931 290605 173959
rect 290639 173931 290667 173959
rect 290701 173931 290729 173959
rect 290763 173931 290791 173959
rect 290577 173869 290605 173897
rect 290639 173869 290667 173897
rect 290701 173869 290729 173897
rect 290763 173869 290791 173897
rect 290577 173807 290605 173835
rect 290639 173807 290667 173835
rect 290701 173807 290729 173835
rect 290763 173807 290791 173835
rect 290577 173745 290605 173773
rect 290639 173745 290667 173773
rect 290701 173745 290729 173773
rect 290763 173745 290791 173773
rect 290577 164931 290605 164959
rect 290639 164931 290667 164959
rect 290701 164931 290729 164959
rect 290763 164931 290791 164959
rect 290577 164869 290605 164897
rect 290639 164869 290667 164897
rect 290701 164869 290729 164897
rect 290763 164869 290791 164897
rect 290577 164807 290605 164835
rect 290639 164807 290667 164835
rect 290701 164807 290729 164835
rect 290763 164807 290791 164835
rect 290577 164745 290605 164773
rect 290639 164745 290667 164773
rect 290701 164745 290729 164773
rect 290763 164745 290791 164773
rect 290577 155931 290605 155959
rect 290639 155931 290667 155959
rect 290701 155931 290729 155959
rect 290763 155931 290791 155959
rect 290577 155869 290605 155897
rect 290639 155869 290667 155897
rect 290701 155869 290729 155897
rect 290763 155869 290791 155897
rect 290577 155807 290605 155835
rect 290639 155807 290667 155835
rect 290701 155807 290729 155835
rect 290763 155807 290791 155835
rect 290577 155745 290605 155773
rect 290639 155745 290667 155773
rect 290701 155745 290729 155773
rect 290763 155745 290791 155773
rect 290577 146931 290605 146959
rect 290639 146931 290667 146959
rect 290701 146931 290729 146959
rect 290763 146931 290791 146959
rect 290577 146869 290605 146897
rect 290639 146869 290667 146897
rect 290701 146869 290729 146897
rect 290763 146869 290791 146897
rect 290577 146807 290605 146835
rect 290639 146807 290667 146835
rect 290701 146807 290729 146835
rect 290763 146807 290791 146835
rect 290577 146745 290605 146773
rect 290639 146745 290667 146773
rect 290701 146745 290729 146773
rect 290763 146745 290791 146773
rect 290577 137931 290605 137959
rect 290639 137931 290667 137959
rect 290701 137931 290729 137959
rect 290763 137931 290791 137959
rect 290577 137869 290605 137897
rect 290639 137869 290667 137897
rect 290701 137869 290729 137897
rect 290763 137869 290791 137897
rect 290577 137807 290605 137835
rect 290639 137807 290667 137835
rect 290701 137807 290729 137835
rect 290763 137807 290791 137835
rect 290577 137745 290605 137773
rect 290639 137745 290667 137773
rect 290701 137745 290729 137773
rect 290763 137745 290791 137773
rect 290577 128931 290605 128959
rect 290639 128931 290667 128959
rect 290701 128931 290729 128959
rect 290763 128931 290791 128959
rect 290577 128869 290605 128897
rect 290639 128869 290667 128897
rect 290701 128869 290729 128897
rect 290763 128869 290791 128897
rect 290577 128807 290605 128835
rect 290639 128807 290667 128835
rect 290701 128807 290729 128835
rect 290763 128807 290791 128835
rect 290577 128745 290605 128773
rect 290639 128745 290667 128773
rect 290701 128745 290729 128773
rect 290763 128745 290791 128773
rect 290577 119931 290605 119959
rect 290639 119931 290667 119959
rect 290701 119931 290729 119959
rect 290763 119931 290791 119959
rect 290577 119869 290605 119897
rect 290639 119869 290667 119897
rect 290701 119869 290729 119897
rect 290763 119869 290791 119897
rect 290577 119807 290605 119835
rect 290639 119807 290667 119835
rect 290701 119807 290729 119835
rect 290763 119807 290791 119835
rect 290577 119745 290605 119773
rect 290639 119745 290667 119773
rect 290701 119745 290729 119773
rect 290763 119745 290791 119773
rect 290577 110931 290605 110959
rect 290639 110931 290667 110959
rect 290701 110931 290729 110959
rect 290763 110931 290791 110959
rect 290577 110869 290605 110897
rect 290639 110869 290667 110897
rect 290701 110869 290729 110897
rect 290763 110869 290791 110897
rect 290577 110807 290605 110835
rect 290639 110807 290667 110835
rect 290701 110807 290729 110835
rect 290763 110807 290791 110835
rect 290577 110745 290605 110773
rect 290639 110745 290667 110773
rect 290701 110745 290729 110773
rect 290763 110745 290791 110773
rect 290577 101931 290605 101959
rect 290639 101931 290667 101959
rect 290701 101931 290729 101959
rect 290763 101931 290791 101959
rect 290577 101869 290605 101897
rect 290639 101869 290667 101897
rect 290701 101869 290729 101897
rect 290763 101869 290791 101897
rect 290577 101807 290605 101835
rect 290639 101807 290667 101835
rect 290701 101807 290729 101835
rect 290763 101807 290791 101835
rect 290577 101745 290605 101773
rect 290639 101745 290667 101773
rect 290701 101745 290729 101773
rect 290763 101745 290791 101773
rect 290577 92931 290605 92959
rect 290639 92931 290667 92959
rect 290701 92931 290729 92959
rect 290763 92931 290791 92959
rect 290577 92869 290605 92897
rect 290639 92869 290667 92897
rect 290701 92869 290729 92897
rect 290763 92869 290791 92897
rect 290577 92807 290605 92835
rect 290639 92807 290667 92835
rect 290701 92807 290729 92835
rect 290763 92807 290791 92835
rect 290577 92745 290605 92773
rect 290639 92745 290667 92773
rect 290701 92745 290729 92773
rect 290763 92745 290791 92773
rect 290577 83931 290605 83959
rect 290639 83931 290667 83959
rect 290701 83931 290729 83959
rect 290763 83931 290791 83959
rect 290577 83869 290605 83897
rect 290639 83869 290667 83897
rect 290701 83869 290729 83897
rect 290763 83869 290791 83897
rect 290577 83807 290605 83835
rect 290639 83807 290667 83835
rect 290701 83807 290729 83835
rect 290763 83807 290791 83835
rect 290577 83745 290605 83773
rect 290639 83745 290667 83773
rect 290701 83745 290729 83773
rect 290763 83745 290791 83773
rect 290577 74931 290605 74959
rect 290639 74931 290667 74959
rect 290701 74931 290729 74959
rect 290763 74931 290791 74959
rect 290577 74869 290605 74897
rect 290639 74869 290667 74897
rect 290701 74869 290729 74897
rect 290763 74869 290791 74897
rect 290577 74807 290605 74835
rect 290639 74807 290667 74835
rect 290701 74807 290729 74835
rect 290763 74807 290791 74835
rect 290577 74745 290605 74773
rect 290639 74745 290667 74773
rect 290701 74745 290729 74773
rect 290763 74745 290791 74773
rect 290577 65931 290605 65959
rect 290639 65931 290667 65959
rect 290701 65931 290729 65959
rect 290763 65931 290791 65959
rect 290577 65869 290605 65897
rect 290639 65869 290667 65897
rect 290701 65869 290729 65897
rect 290763 65869 290791 65897
rect 290577 65807 290605 65835
rect 290639 65807 290667 65835
rect 290701 65807 290729 65835
rect 290763 65807 290791 65835
rect 290577 65745 290605 65773
rect 290639 65745 290667 65773
rect 290701 65745 290729 65773
rect 290763 65745 290791 65773
rect 290577 56931 290605 56959
rect 290639 56931 290667 56959
rect 290701 56931 290729 56959
rect 290763 56931 290791 56959
rect 290577 56869 290605 56897
rect 290639 56869 290667 56897
rect 290701 56869 290729 56897
rect 290763 56869 290791 56897
rect 290577 56807 290605 56835
rect 290639 56807 290667 56835
rect 290701 56807 290729 56835
rect 290763 56807 290791 56835
rect 290577 56745 290605 56773
rect 290639 56745 290667 56773
rect 290701 56745 290729 56773
rect 290763 56745 290791 56773
rect 290577 47931 290605 47959
rect 290639 47931 290667 47959
rect 290701 47931 290729 47959
rect 290763 47931 290791 47959
rect 290577 47869 290605 47897
rect 290639 47869 290667 47897
rect 290701 47869 290729 47897
rect 290763 47869 290791 47897
rect 290577 47807 290605 47835
rect 290639 47807 290667 47835
rect 290701 47807 290729 47835
rect 290763 47807 290791 47835
rect 290577 47745 290605 47773
rect 290639 47745 290667 47773
rect 290701 47745 290729 47773
rect 290763 47745 290791 47773
rect 290577 38931 290605 38959
rect 290639 38931 290667 38959
rect 290701 38931 290729 38959
rect 290763 38931 290791 38959
rect 290577 38869 290605 38897
rect 290639 38869 290667 38897
rect 290701 38869 290729 38897
rect 290763 38869 290791 38897
rect 290577 38807 290605 38835
rect 290639 38807 290667 38835
rect 290701 38807 290729 38835
rect 290763 38807 290791 38835
rect 290577 38745 290605 38773
rect 290639 38745 290667 38773
rect 290701 38745 290729 38773
rect 290763 38745 290791 38773
rect 290577 29931 290605 29959
rect 290639 29931 290667 29959
rect 290701 29931 290729 29959
rect 290763 29931 290791 29959
rect 290577 29869 290605 29897
rect 290639 29869 290667 29897
rect 290701 29869 290729 29897
rect 290763 29869 290791 29897
rect 290577 29807 290605 29835
rect 290639 29807 290667 29835
rect 290701 29807 290729 29835
rect 290763 29807 290791 29835
rect 290577 29745 290605 29773
rect 290639 29745 290667 29773
rect 290701 29745 290729 29773
rect 290763 29745 290791 29773
rect 290577 20931 290605 20959
rect 290639 20931 290667 20959
rect 290701 20931 290729 20959
rect 290763 20931 290791 20959
rect 290577 20869 290605 20897
rect 290639 20869 290667 20897
rect 290701 20869 290729 20897
rect 290763 20869 290791 20897
rect 290577 20807 290605 20835
rect 290639 20807 290667 20835
rect 290701 20807 290729 20835
rect 290763 20807 290791 20835
rect 290577 20745 290605 20773
rect 290639 20745 290667 20773
rect 290701 20745 290729 20773
rect 290763 20745 290791 20773
rect 290577 11931 290605 11959
rect 290639 11931 290667 11959
rect 290701 11931 290729 11959
rect 290763 11931 290791 11959
rect 290577 11869 290605 11897
rect 290639 11869 290667 11897
rect 290701 11869 290729 11897
rect 290763 11869 290791 11897
rect 290577 11807 290605 11835
rect 290639 11807 290667 11835
rect 290701 11807 290729 11835
rect 290763 11807 290791 11835
rect 290577 11745 290605 11773
rect 290639 11745 290667 11773
rect 290701 11745 290729 11773
rect 290763 11745 290791 11773
rect 290577 2931 290605 2959
rect 290639 2931 290667 2959
rect 290701 2931 290729 2959
rect 290763 2931 290791 2959
rect 290577 2869 290605 2897
rect 290639 2869 290667 2897
rect 290701 2869 290729 2897
rect 290763 2869 290791 2897
rect 290577 2807 290605 2835
rect 290639 2807 290667 2835
rect 290701 2807 290729 2835
rect 290763 2807 290791 2835
rect 290577 2745 290605 2773
rect 290639 2745 290667 2773
rect 290701 2745 290729 2773
rect 290763 2745 290791 2773
rect 290577 876 290605 904
rect 290639 876 290667 904
rect 290701 876 290729 904
rect 290763 876 290791 904
rect 290577 814 290605 842
rect 290639 814 290667 842
rect 290701 814 290729 842
rect 290763 814 290791 842
rect 290577 752 290605 780
rect 290639 752 290667 780
rect 290701 752 290729 780
rect 290763 752 290791 780
rect 290577 690 290605 718
rect 290639 690 290667 718
rect 290701 690 290729 718
rect 290763 690 290791 718
rect 292437 299642 292465 299670
rect 292499 299642 292527 299670
rect 292561 299642 292589 299670
rect 292623 299642 292651 299670
rect 292437 299580 292465 299608
rect 292499 299580 292527 299608
rect 292561 299580 292589 299608
rect 292623 299580 292651 299608
rect 292437 299518 292465 299546
rect 292499 299518 292527 299546
rect 292561 299518 292589 299546
rect 292623 299518 292651 299546
rect 292437 299456 292465 299484
rect 292499 299456 292527 299484
rect 292561 299456 292589 299484
rect 292623 299456 292651 299484
rect 299736 299642 299764 299670
rect 299798 299642 299826 299670
rect 299860 299642 299888 299670
rect 299922 299642 299950 299670
rect 299736 299580 299764 299608
rect 299798 299580 299826 299608
rect 299860 299580 299888 299608
rect 299922 299580 299950 299608
rect 299736 299518 299764 299546
rect 299798 299518 299826 299546
rect 299860 299518 299888 299546
rect 299922 299518 299950 299546
rect 299736 299456 299764 299484
rect 299798 299456 299826 299484
rect 299860 299456 299888 299484
rect 299922 299456 299950 299484
rect 292437 293931 292465 293959
rect 292499 293931 292527 293959
rect 292561 293931 292589 293959
rect 292623 293931 292651 293959
rect 292437 293869 292465 293897
rect 292499 293869 292527 293897
rect 292561 293869 292589 293897
rect 292623 293869 292651 293897
rect 292437 293807 292465 293835
rect 292499 293807 292527 293835
rect 292561 293807 292589 293835
rect 292623 293807 292651 293835
rect 292437 293745 292465 293773
rect 292499 293745 292527 293773
rect 292561 293745 292589 293773
rect 292623 293745 292651 293773
rect 292437 284931 292465 284959
rect 292499 284931 292527 284959
rect 292561 284931 292589 284959
rect 292623 284931 292651 284959
rect 292437 284869 292465 284897
rect 292499 284869 292527 284897
rect 292561 284869 292589 284897
rect 292623 284869 292651 284897
rect 292437 284807 292465 284835
rect 292499 284807 292527 284835
rect 292561 284807 292589 284835
rect 292623 284807 292651 284835
rect 292437 284745 292465 284773
rect 292499 284745 292527 284773
rect 292561 284745 292589 284773
rect 292623 284745 292651 284773
rect 292437 275931 292465 275959
rect 292499 275931 292527 275959
rect 292561 275931 292589 275959
rect 292623 275931 292651 275959
rect 292437 275869 292465 275897
rect 292499 275869 292527 275897
rect 292561 275869 292589 275897
rect 292623 275869 292651 275897
rect 292437 275807 292465 275835
rect 292499 275807 292527 275835
rect 292561 275807 292589 275835
rect 292623 275807 292651 275835
rect 292437 275745 292465 275773
rect 292499 275745 292527 275773
rect 292561 275745 292589 275773
rect 292623 275745 292651 275773
rect 292437 266931 292465 266959
rect 292499 266931 292527 266959
rect 292561 266931 292589 266959
rect 292623 266931 292651 266959
rect 292437 266869 292465 266897
rect 292499 266869 292527 266897
rect 292561 266869 292589 266897
rect 292623 266869 292651 266897
rect 292437 266807 292465 266835
rect 292499 266807 292527 266835
rect 292561 266807 292589 266835
rect 292623 266807 292651 266835
rect 292437 266745 292465 266773
rect 292499 266745 292527 266773
rect 292561 266745 292589 266773
rect 292623 266745 292651 266773
rect 292437 257931 292465 257959
rect 292499 257931 292527 257959
rect 292561 257931 292589 257959
rect 292623 257931 292651 257959
rect 292437 257869 292465 257897
rect 292499 257869 292527 257897
rect 292561 257869 292589 257897
rect 292623 257869 292651 257897
rect 292437 257807 292465 257835
rect 292499 257807 292527 257835
rect 292561 257807 292589 257835
rect 292623 257807 292651 257835
rect 292437 257745 292465 257773
rect 292499 257745 292527 257773
rect 292561 257745 292589 257773
rect 292623 257745 292651 257773
rect 292437 248931 292465 248959
rect 292499 248931 292527 248959
rect 292561 248931 292589 248959
rect 292623 248931 292651 248959
rect 292437 248869 292465 248897
rect 292499 248869 292527 248897
rect 292561 248869 292589 248897
rect 292623 248869 292651 248897
rect 292437 248807 292465 248835
rect 292499 248807 292527 248835
rect 292561 248807 292589 248835
rect 292623 248807 292651 248835
rect 292437 248745 292465 248773
rect 292499 248745 292527 248773
rect 292561 248745 292589 248773
rect 292623 248745 292651 248773
rect 292437 239931 292465 239959
rect 292499 239931 292527 239959
rect 292561 239931 292589 239959
rect 292623 239931 292651 239959
rect 292437 239869 292465 239897
rect 292499 239869 292527 239897
rect 292561 239869 292589 239897
rect 292623 239869 292651 239897
rect 292437 239807 292465 239835
rect 292499 239807 292527 239835
rect 292561 239807 292589 239835
rect 292623 239807 292651 239835
rect 292437 239745 292465 239773
rect 292499 239745 292527 239773
rect 292561 239745 292589 239773
rect 292623 239745 292651 239773
rect 292437 230931 292465 230959
rect 292499 230931 292527 230959
rect 292561 230931 292589 230959
rect 292623 230931 292651 230959
rect 292437 230869 292465 230897
rect 292499 230869 292527 230897
rect 292561 230869 292589 230897
rect 292623 230869 292651 230897
rect 292437 230807 292465 230835
rect 292499 230807 292527 230835
rect 292561 230807 292589 230835
rect 292623 230807 292651 230835
rect 292437 230745 292465 230773
rect 292499 230745 292527 230773
rect 292561 230745 292589 230773
rect 292623 230745 292651 230773
rect 292437 221931 292465 221959
rect 292499 221931 292527 221959
rect 292561 221931 292589 221959
rect 292623 221931 292651 221959
rect 292437 221869 292465 221897
rect 292499 221869 292527 221897
rect 292561 221869 292589 221897
rect 292623 221869 292651 221897
rect 292437 221807 292465 221835
rect 292499 221807 292527 221835
rect 292561 221807 292589 221835
rect 292623 221807 292651 221835
rect 292437 221745 292465 221773
rect 292499 221745 292527 221773
rect 292561 221745 292589 221773
rect 292623 221745 292651 221773
rect 292437 212931 292465 212959
rect 292499 212931 292527 212959
rect 292561 212931 292589 212959
rect 292623 212931 292651 212959
rect 292437 212869 292465 212897
rect 292499 212869 292527 212897
rect 292561 212869 292589 212897
rect 292623 212869 292651 212897
rect 292437 212807 292465 212835
rect 292499 212807 292527 212835
rect 292561 212807 292589 212835
rect 292623 212807 292651 212835
rect 292437 212745 292465 212773
rect 292499 212745 292527 212773
rect 292561 212745 292589 212773
rect 292623 212745 292651 212773
rect 292437 203931 292465 203959
rect 292499 203931 292527 203959
rect 292561 203931 292589 203959
rect 292623 203931 292651 203959
rect 292437 203869 292465 203897
rect 292499 203869 292527 203897
rect 292561 203869 292589 203897
rect 292623 203869 292651 203897
rect 292437 203807 292465 203835
rect 292499 203807 292527 203835
rect 292561 203807 292589 203835
rect 292623 203807 292651 203835
rect 292437 203745 292465 203773
rect 292499 203745 292527 203773
rect 292561 203745 292589 203773
rect 292623 203745 292651 203773
rect 292437 194931 292465 194959
rect 292499 194931 292527 194959
rect 292561 194931 292589 194959
rect 292623 194931 292651 194959
rect 292437 194869 292465 194897
rect 292499 194869 292527 194897
rect 292561 194869 292589 194897
rect 292623 194869 292651 194897
rect 292437 194807 292465 194835
rect 292499 194807 292527 194835
rect 292561 194807 292589 194835
rect 292623 194807 292651 194835
rect 292437 194745 292465 194773
rect 292499 194745 292527 194773
rect 292561 194745 292589 194773
rect 292623 194745 292651 194773
rect 292437 185931 292465 185959
rect 292499 185931 292527 185959
rect 292561 185931 292589 185959
rect 292623 185931 292651 185959
rect 292437 185869 292465 185897
rect 292499 185869 292527 185897
rect 292561 185869 292589 185897
rect 292623 185869 292651 185897
rect 292437 185807 292465 185835
rect 292499 185807 292527 185835
rect 292561 185807 292589 185835
rect 292623 185807 292651 185835
rect 292437 185745 292465 185773
rect 292499 185745 292527 185773
rect 292561 185745 292589 185773
rect 292623 185745 292651 185773
rect 292437 176931 292465 176959
rect 292499 176931 292527 176959
rect 292561 176931 292589 176959
rect 292623 176931 292651 176959
rect 292437 176869 292465 176897
rect 292499 176869 292527 176897
rect 292561 176869 292589 176897
rect 292623 176869 292651 176897
rect 292437 176807 292465 176835
rect 292499 176807 292527 176835
rect 292561 176807 292589 176835
rect 292623 176807 292651 176835
rect 292437 176745 292465 176773
rect 292499 176745 292527 176773
rect 292561 176745 292589 176773
rect 292623 176745 292651 176773
rect 292437 167931 292465 167959
rect 292499 167931 292527 167959
rect 292561 167931 292589 167959
rect 292623 167931 292651 167959
rect 292437 167869 292465 167897
rect 292499 167869 292527 167897
rect 292561 167869 292589 167897
rect 292623 167869 292651 167897
rect 292437 167807 292465 167835
rect 292499 167807 292527 167835
rect 292561 167807 292589 167835
rect 292623 167807 292651 167835
rect 292437 167745 292465 167773
rect 292499 167745 292527 167773
rect 292561 167745 292589 167773
rect 292623 167745 292651 167773
rect 292437 158931 292465 158959
rect 292499 158931 292527 158959
rect 292561 158931 292589 158959
rect 292623 158931 292651 158959
rect 292437 158869 292465 158897
rect 292499 158869 292527 158897
rect 292561 158869 292589 158897
rect 292623 158869 292651 158897
rect 292437 158807 292465 158835
rect 292499 158807 292527 158835
rect 292561 158807 292589 158835
rect 292623 158807 292651 158835
rect 292437 158745 292465 158773
rect 292499 158745 292527 158773
rect 292561 158745 292589 158773
rect 292623 158745 292651 158773
rect 292437 149931 292465 149959
rect 292499 149931 292527 149959
rect 292561 149931 292589 149959
rect 292623 149931 292651 149959
rect 292437 149869 292465 149897
rect 292499 149869 292527 149897
rect 292561 149869 292589 149897
rect 292623 149869 292651 149897
rect 292437 149807 292465 149835
rect 292499 149807 292527 149835
rect 292561 149807 292589 149835
rect 292623 149807 292651 149835
rect 292437 149745 292465 149773
rect 292499 149745 292527 149773
rect 292561 149745 292589 149773
rect 292623 149745 292651 149773
rect 292437 140931 292465 140959
rect 292499 140931 292527 140959
rect 292561 140931 292589 140959
rect 292623 140931 292651 140959
rect 292437 140869 292465 140897
rect 292499 140869 292527 140897
rect 292561 140869 292589 140897
rect 292623 140869 292651 140897
rect 292437 140807 292465 140835
rect 292499 140807 292527 140835
rect 292561 140807 292589 140835
rect 292623 140807 292651 140835
rect 292437 140745 292465 140773
rect 292499 140745 292527 140773
rect 292561 140745 292589 140773
rect 292623 140745 292651 140773
rect 292437 131931 292465 131959
rect 292499 131931 292527 131959
rect 292561 131931 292589 131959
rect 292623 131931 292651 131959
rect 292437 131869 292465 131897
rect 292499 131869 292527 131897
rect 292561 131869 292589 131897
rect 292623 131869 292651 131897
rect 292437 131807 292465 131835
rect 292499 131807 292527 131835
rect 292561 131807 292589 131835
rect 292623 131807 292651 131835
rect 292437 131745 292465 131773
rect 292499 131745 292527 131773
rect 292561 131745 292589 131773
rect 292623 131745 292651 131773
rect 292437 122931 292465 122959
rect 292499 122931 292527 122959
rect 292561 122931 292589 122959
rect 292623 122931 292651 122959
rect 292437 122869 292465 122897
rect 292499 122869 292527 122897
rect 292561 122869 292589 122897
rect 292623 122869 292651 122897
rect 292437 122807 292465 122835
rect 292499 122807 292527 122835
rect 292561 122807 292589 122835
rect 292623 122807 292651 122835
rect 292437 122745 292465 122773
rect 292499 122745 292527 122773
rect 292561 122745 292589 122773
rect 292623 122745 292651 122773
rect 292437 113931 292465 113959
rect 292499 113931 292527 113959
rect 292561 113931 292589 113959
rect 292623 113931 292651 113959
rect 292437 113869 292465 113897
rect 292499 113869 292527 113897
rect 292561 113869 292589 113897
rect 292623 113869 292651 113897
rect 292437 113807 292465 113835
rect 292499 113807 292527 113835
rect 292561 113807 292589 113835
rect 292623 113807 292651 113835
rect 292437 113745 292465 113773
rect 292499 113745 292527 113773
rect 292561 113745 292589 113773
rect 292623 113745 292651 113773
rect 292437 104931 292465 104959
rect 292499 104931 292527 104959
rect 292561 104931 292589 104959
rect 292623 104931 292651 104959
rect 292437 104869 292465 104897
rect 292499 104869 292527 104897
rect 292561 104869 292589 104897
rect 292623 104869 292651 104897
rect 292437 104807 292465 104835
rect 292499 104807 292527 104835
rect 292561 104807 292589 104835
rect 292623 104807 292651 104835
rect 292437 104745 292465 104773
rect 292499 104745 292527 104773
rect 292561 104745 292589 104773
rect 292623 104745 292651 104773
rect 292437 95931 292465 95959
rect 292499 95931 292527 95959
rect 292561 95931 292589 95959
rect 292623 95931 292651 95959
rect 292437 95869 292465 95897
rect 292499 95869 292527 95897
rect 292561 95869 292589 95897
rect 292623 95869 292651 95897
rect 292437 95807 292465 95835
rect 292499 95807 292527 95835
rect 292561 95807 292589 95835
rect 292623 95807 292651 95835
rect 292437 95745 292465 95773
rect 292499 95745 292527 95773
rect 292561 95745 292589 95773
rect 292623 95745 292651 95773
rect 292437 86931 292465 86959
rect 292499 86931 292527 86959
rect 292561 86931 292589 86959
rect 292623 86931 292651 86959
rect 292437 86869 292465 86897
rect 292499 86869 292527 86897
rect 292561 86869 292589 86897
rect 292623 86869 292651 86897
rect 292437 86807 292465 86835
rect 292499 86807 292527 86835
rect 292561 86807 292589 86835
rect 292623 86807 292651 86835
rect 292437 86745 292465 86773
rect 292499 86745 292527 86773
rect 292561 86745 292589 86773
rect 292623 86745 292651 86773
rect 292437 77931 292465 77959
rect 292499 77931 292527 77959
rect 292561 77931 292589 77959
rect 292623 77931 292651 77959
rect 292437 77869 292465 77897
rect 292499 77869 292527 77897
rect 292561 77869 292589 77897
rect 292623 77869 292651 77897
rect 292437 77807 292465 77835
rect 292499 77807 292527 77835
rect 292561 77807 292589 77835
rect 292623 77807 292651 77835
rect 292437 77745 292465 77773
rect 292499 77745 292527 77773
rect 292561 77745 292589 77773
rect 292623 77745 292651 77773
rect 292437 68931 292465 68959
rect 292499 68931 292527 68959
rect 292561 68931 292589 68959
rect 292623 68931 292651 68959
rect 292437 68869 292465 68897
rect 292499 68869 292527 68897
rect 292561 68869 292589 68897
rect 292623 68869 292651 68897
rect 292437 68807 292465 68835
rect 292499 68807 292527 68835
rect 292561 68807 292589 68835
rect 292623 68807 292651 68835
rect 292437 68745 292465 68773
rect 292499 68745 292527 68773
rect 292561 68745 292589 68773
rect 292623 68745 292651 68773
rect 292437 59931 292465 59959
rect 292499 59931 292527 59959
rect 292561 59931 292589 59959
rect 292623 59931 292651 59959
rect 292437 59869 292465 59897
rect 292499 59869 292527 59897
rect 292561 59869 292589 59897
rect 292623 59869 292651 59897
rect 292437 59807 292465 59835
rect 292499 59807 292527 59835
rect 292561 59807 292589 59835
rect 292623 59807 292651 59835
rect 292437 59745 292465 59773
rect 292499 59745 292527 59773
rect 292561 59745 292589 59773
rect 292623 59745 292651 59773
rect 292437 50931 292465 50959
rect 292499 50931 292527 50959
rect 292561 50931 292589 50959
rect 292623 50931 292651 50959
rect 292437 50869 292465 50897
rect 292499 50869 292527 50897
rect 292561 50869 292589 50897
rect 292623 50869 292651 50897
rect 292437 50807 292465 50835
rect 292499 50807 292527 50835
rect 292561 50807 292589 50835
rect 292623 50807 292651 50835
rect 292437 50745 292465 50773
rect 292499 50745 292527 50773
rect 292561 50745 292589 50773
rect 292623 50745 292651 50773
rect 292437 41931 292465 41959
rect 292499 41931 292527 41959
rect 292561 41931 292589 41959
rect 292623 41931 292651 41959
rect 292437 41869 292465 41897
rect 292499 41869 292527 41897
rect 292561 41869 292589 41897
rect 292623 41869 292651 41897
rect 292437 41807 292465 41835
rect 292499 41807 292527 41835
rect 292561 41807 292589 41835
rect 292623 41807 292651 41835
rect 292437 41745 292465 41773
rect 292499 41745 292527 41773
rect 292561 41745 292589 41773
rect 292623 41745 292651 41773
rect 292437 32931 292465 32959
rect 292499 32931 292527 32959
rect 292561 32931 292589 32959
rect 292623 32931 292651 32959
rect 292437 32869 292465 32897
rect 292499 32869 292527 32897
rect 292561 32869 292589 32897
rect 292623 32869 292651 32897
rect 292437 32807 292465 32835
rect 292499 32807 292527 32835
rect 292561 32807 292589 32835
rect 292623 32807 292651 32835
rect 292437 32745 292465 32773
rect 292499 32745 292527 32773
rect 292561 32745 292589 32773
rect 292623 32745 292651 32773
rect 292437 23931 292465 23959
rect 292499 23931 292527 23959
rect 292561 23931 292589 23959
rect 292623 23931 292651 23959
rect 292437 23869 292465 23897
rect 292499 23869 292527 23897
rect 292561 23869 292589 23897
rect 292623 23869 292651 23897
rect 292437 23807 292465 23835
rect 292499 23807 292527 23835
rect 292561 23807 292589 23835
rect 292623 23807 292651 23835
rect 292437 23745 292465 23773
rect 292499 23745 292527 23773
rect 292561 23745 292589 23773
rect 292623 23745 292651 23773
rect 292437 14931 292465 14959
rect 292499 14931 292527 14959
rect 292561 14931 292589 14959
rect 292623 14931 292651 14959
rect 292437 14869 292465 14897
rect 292499 14869 292527 14897
rect 292561 14869 292589 14897
rect 292623 14869 292651 14897
rect 292437 14807 292465 14835
rect 292499 14807 292527 14835
rect 292561 14807 292589 14835
rect 292623 14807 292651 14835
rect 292437 14745 292465 14773
rect 292499 14745 292527 14773
rect 292561 14745 292589 14773
rect 292623 14745 292651 14773
rect 292437 5931 292465 5959
rect 292499 5931 292527 5959
rect 292561 5931 292589 5959
rect 292623 5931 292651 5959
rect 292437 5869 292465 5897
rect 292499 5869 292527 5897
rect 292561 5869 292589 5897
rect 292623 5869 292651 5897
rect 292437 5807 292465 5835
rect 292499 5807 292527 5835
rect 292561 5807 292589 5835
rect 292623 5807 292651 5835
rect 292437 5745 292465 5773
rect 292499 5745 292527 5773
rect 292561 5745 292589 5773
rect 292623 5745 292651 5773
rect 299256 299162 299284 299190
rect 299318 299162 299346 299190
rect 299380 299162 299408 299190
rect 299442 299162 299470 299190
rect 299256 299100 299284 299128
rect 299318 299100 299346 299128
rect 299380 299100 299408 299128
rect 299442 299100 299470 299128
rect 299256 299038 299284 299066
rect 299318 299038 299346 299066
rect 299380 299038 299408 299066
rect 299442 299038 299470 299066
rect 299256 298976 299284 299004
rect 299318 298976 299346 299004
rect 299380 298976 299408 299004
rect 299442 298976 299470 299004
rect 299256 290931 299284 290959
rect 299318 290931 299346 290959
rect 299380 290931 299408 290959
rect 299442 290931 299470 290959
rect 299256 290869 299284 290897
rect 299318 290869 299346 290897
rect 299380 290869 299408 290897
rect 299442 290869 299470 290897
rect 299256 290807 299284 290835
rect 299318 290807 299346 290835
rect 299380 290807 299408 290835
rect 299442 290807 299470 290835
rect 299256 290745 299284 290773
rect 299318 290745 299346 290773
rect 299380 290745 299408 290773
rect 299442 290745 299470 290773
rect 299256 281931 299284 281959
rect 299318 281931 299346 281959
rect 299380 281931 299408 281959
rect 299442 281931 299470 281959
rect 299256 281869 299284 281897
rect 299318 281869 299346 281897
rect 299380 281869 299408 281897
rect 299442 281869 299470 281897
rect 299256 281807 299284 281835
rect 299318 281807 299346 281835
rect 299380 281807 299408 281835
rect 299442 281807 299470 281835
rect 299256 281745 299284 281773
rect 299318 281745 299346 281773
rect 299380 281745 299408 281773
rect 299442 281745 299470 281773
rect 299256 272931 299284 272959
rect 299318 272931 299346 272959
rect 299380 272931 299408 272959
rect 299442 272931 299470 272959
rect 299256 272869 299284 272897
rect 299318 272869 299346 272897
rect 299380 272869 299408 272897
rect 299442 272869 299470 272897
rect 299256 272807 299284 272835
rect 299318 272807 299346 272835
rect 299380 272807 299408 272835
rect 299442 272807 299470 272835
rect 299256 272745 299284 272773
rect 299318 272745 299346 272773
rect 299380 272745 299408 272773
rect 299442 272745 299470 272773
rect 299256 263931 299284 263959
rect 299318 263931 299346 263959
rect 299380 263931 299408 263959
rect 299442 263931 299470 263959
rect 299256 263869 299284 263897
rect 299318 263869 299346 263897
rect 299380 263869 299408 263897
rect 299442 263869 299470 263897
rect 299256 263807 299284 263835
rect 299318 263807 299346 263835
rect 299380 263807 299408 263835
rect 299442 263807 299470 263835
rect 299256 263745 299284 263773
rect 299318 263745 299346 263773
rect 299380 263745 299408 263773
rect 299442 263745 299470 263773
rect 299256 254931 299284 254959
rect 299318 254931 299346 254959
rect 299380 254931 299408 254959
rect 299442 254931 299470 254959
rect 299256 254869 299284 254897
rect 299318 254869 299346 254897
rect 299380 254869 299408 254897
rect 299442 254869 299470 254897
rect 299256 254807 299284 254835
rect 299318 254807 299346 254835
rect 299380 254807 299408 254835
rect 299442 254807 299470 254835
rect 299256 254745 299284 254773
rect 299318 254745 299346 254773
rect 299380 254745 299408 254773
rect 299442 254745 299470 254773
rect 299256 245931 299284 245959
rect 299318 245931 299346 245959
rect 299380 245931 299408 245959
rect 299442 245931 299470 245959
rect 299256 245869 299284 245897
rect 299318 245869 299346 245897
rect 299380 245869 299408 245897
rect 299442 245869 299470 245897
rect 299256 245807 299284 245835
rect 299318 245807 299346 245835
rect 299380 245807 299408 245835
rect 299442 245807 299470 245835
rect 299256 245745 299284 245773
rect 299318 245745 299346 245773
rect 299380 245745 299408 245773
rect 299442 245745 299470 245773
rect 299256 236931 299284 236959
rect 299318 236931 299346 236959
rect 299380 236931 299408 236959
rect 299442 236931 299470 236959
rect 299256 236869 299284 236897
rect 299318 236869 299346 236897
rect 299380 236869 299408 236897
rect 299442 236869 299470 236897
rect 299256 236807 299284 236835
rect 299318 236807 299346 236835
rect 299380 236807 299408 236835
rect 299442 236807 299470 236835
rect 299256 236745 299284 236773
rect 299318 236745 299346 236773
rect 299380 236745 299408 236773
rect 299442 236745 299470 236773
rect 299256 227931 299284 227959
rect 299318 227931 299346 227959
rect 299380 227931 299408 227959
rect 299442 227931 299470 227959
rect 299256 227869 299284 227897
rect 299318 227869 299346 227897
rect 299380 227869 299408 227897
rect 299442 227869 299470 227897
rect 299256 227807 299284 227835
rect 299318 227807 299346 227835
rect 299380 227807 299408 227835
rect 299442 227807 299470 227835
rect 299256 227745 299284 227773
rect 299318 227745 299346 227773
rect 299380 227745 299408 227773
rect 299442 227745 299470 227773
rect 299256 218931 299284 218959
rect 299318 218931 299346 218959
rect 299380 218931 299408 218959
rect 299442 218931 299470 218959
rect 299256 218869 299284 218897
rect 299318 218869 299346 218897
rect 299380 218869 299408 218897
rect 299442 218869 299470 218897
rect 299256 218807 299284 218835
rect 299318 218807 299346 218835
rect 299380 218807 299408 218835
rect 299442 218807 299470 218835
rect 299256 218745 299284 218773
rect 299318 218745 299346 218773
rect 299380 218745 299408 218773
rect 299442 218745 299470 218773
rect 299256 209931 299284 209959
rect 299318 209931 299346 209959
rect 299380 209931 299408 209959
rect 299442 209931 299470 209959
rect 299256 209869 299284 209897
rect 299318 209869 299346 209897
rect 299380 209869 299408 209897
rect 299442 209869 299470 209897
rect 299256 209807 299284 209835
rect 299318 209807 299346 209835
rect 299380 209807 299408 209835
rect 299442 209807 299470 209835
rect 299256 209745 299284 209773
rect 299318 209745 299346 209773
rect 299380 209745 299408 209773
rect 299442 209745 299470 209773
rect 299256 200931 299284 200959
rect 299318 200931 299346 200959
rect 299380 200931 299408 200959
rect 299442 200931 299470 200959
rect 299256 200869 299284 200897
rect 299318 200869 299346 200897
rect 299380 200869 299408 200897
rect 299442 200869 299470 200897
rect 299256 200807 299284 200835
rect 299318 200807 299346 200835
rect 299380 200807 299408 200835
rect 299442 200807 299470 200835
rect 299256 200745 299284 200773
rect 299318 200745 299346 200773
rect 299380 200745 299408 200773
rect 299442 200745 299470 200773
rect 299256 191931 299284 191959
rect 299318 191931 299346 191959
rect 299380 191931 299408 191959
rect 299442 191931 299470 191959
rect 299256 191869 299284 191897
rect 299318 191869 299346 191897
rect 299380 191869 299408 191897
rect 299442 191869 299470 191897
rect 299256 191807 299284 191835
rect 299318 191807 299346 191835
rect 299380 191807 299408 191835
rect 299442 191807 299470 191835
rect 299256 191745 299284 191773
rect 299318 191745 299346 191773
rect 299380 191745 299408 191773
rect 299442 191745 299470 191773
rect 299256 182931 299284 182959
rect 299318 182931 299346 182959
rect 299380 182931 299408 182959
rect 299442 182931 299470 182959
rect 299256 182869 299284 182897
rect 299318 182869 299346 182897
rect 299380 182869 299408 182897
rect 299442 182869 299470 182897
rect 299256 182807 299284 182835
rect 299318 182807 299346 182835
rect 299380 182807 299408 182835
rect 299442 182807 299470 182835
rect 299256 182745 299284 182773
rect 299318 182745 299346 182773
rect 299380 182745 299408 182773
rect 299442 182745 299470 182773
rect 299256 173931 299284 173959
rect 299318 173931 299346 173959
rect 299380 173931 299408 173959
rect 299442 173931 299470 173959
rect 299256 173869 299284 173897
rect 299318 173869 299346 173897
rect 299380 173869 299408 173897
rect 299442 173869 299470 173897
rect 299256 173807 299284 173835
rect 299318 173807 299346 173835
rect 299380 173807 299408 173835
rect 299442 173807 299470 173835
rect 299256 173745 299284 173773
rect 299318 173745 299346 173773
rect 299380 173745 299408 173773
rect 299442 173745 299470 173773
rect 299256 164931 299284 164959
rect 299318 164931 299346 164959
rect 299380 164931 299408 164959
rect 299442 164931 299470 164959
rect 299256 164869 299284 164897
rect 299318 164869 299346 164897
rect 299380 164869 299408 164897
rect 299442 164869 299470 164897
rect 299256 164807 299284 164835
rect 299318 164807 299346 164835
rect 299380 164807 299408 164835
rect 299442 164807 299470 164835
rect 299256 164745 299284 164773
rect 299318 164745 299346 164773
rect 299380 164745 299408 164773
rect 299442 164745 299470 164773
rect 299256 155931 299284 155959
rect 299318 155931 299346 155959
rect 299380 155931 299408 155959
rect 299442 155931 299470 155959
rect 299256 155869 299284 155897
rect 299318 155869 299346 155897
rect 299380 155869 299408 155897
rect 299442 155869 299470 155897
rect 299256 155807 299284 155835
rect 299318 155807 299346 155835
rect 299380 155807 299408 155835
rect 299442 155807 299470 155835
rect 299256 155745 299284 155773
rect 299318 155745 299346 155773
rect 299380 155745 299408 155773
rect 299442 155745 299470 155773
rect 299256 146931 299284 146959
rect 299318 146931 299346 146959
rect 299380 146931 299408 146959
rect 299442 146931 299470 146959
rect 299256 146869 299284 146897
rect 299318 146869 299346 146897
rect 299380 146869 299408 146897
rect 299442 146869 299470 146897
rect 299256 146807 299284 146835
rect 299318 146807 299346 146835
rect 299380 146807 299408 146835
rect 299442 146807 299470 146835
rect 299256 146745 299284 146773
rect 299318 146745 299346 146773
rect 299380 146745 299408 146773
rect 299442 146745 299470 146773
rect 299256 137931 299284 137959
rect 299318 137931 299346 137959
rect 299380 137931 299408 137959
rect 299442 137931 299470 137959
rect 299256 137869 299284 137897
rect 299318 137869 299346 137897
rect 299380 137869 299408 137897
rect 299442 137869 299470 137897
rect 299256 137807 299284 137835
rect 299318 137807 299346 137835
rect 299380 137807 299408 137835
rect 299442 137807 299470 137835
rect 299256 137745 299284 137773
rect 299318 137745 299346 137773
rect 299380 137745 299408 137773
rect 299442 137745 299470 137773
rect 299256 128931 299284 128959
rect 299318 128931 299346 128959
rect 299380 128931 299408 128959
rect 299442 128931 299470 128959
rect 299256 128869 299284 128897
rect 299318 128869 299346 128897
rect 299380 128869 299408 128897
rect 299442 128869 299470 128897
rect 299256 128807 299284 128835
rect 299318 128807 299346 128835
rect 299380 128807 299408 128835
rect 299442 128807 299470 128835
rect 299256 128745 299284 128773
rect 299318 128745 299346 128773
rect 299380 128745 299408 128773
rect 299442 128745 299470 128773
rect 299256 119931 299284 119959
rect 299318 119931 299346 119959
rect 299380 119931 299408 119959
rect 299442 119931 299470 119959
rect 299256 119869 299284 119897
rect 299318 119869 299346 119897
rect 299380 119869 299408 119897
rect 299442 119869 299470 119897
rect 299256 119807 299284 119835
rect 299318 119807 299346 119835
rect 299380 119807 299408 119835
rect 299442 119807 299470 119835
rect 299256 119745 299284 119773
rect 299318 119745 299346 119773
rect 299380 119745 299408 119773
rect 299442 119745 299470 119773
rect 299256 110931 299284 110959
rect 299318 110931 299346 110959
rect 299380 110931 299408 110959
rect 299442 110931 299470 110959
rect 299256 110869 299284 110897
rect 299318 110869 299346 110897
rect 299380 110869 299408 110897
rect 299442 110869 299470 110897
rect 299256 110807 299284 110835
rect 299318 110807 299346 110835
rect 299380 110807 299408 110835
rect 299442 110807 299470 110835
rect 299256 110745 299284 110773
rect 299318 110745 299346 110773
rect 299380 110745 299408 110773
rect 299442 110745 299470 110773
rect 299256 101931 299284 101959
rect 299318 101931 299346 101959
rect 299380 101931 299408 101959
rect 299442 101931 299470 101959
rect 299256 101869 299284 101897
rect 299318 101869 299346 101897
rect 299380 101869 299408 101897
rect 299442 101869 299470 101897
rect 299256 101807 299284 101835
rect 299318 101807 299346 101835
rect 299380 101807 299408 101835
rect 299442 101807 299470 101835
rect 299256 101745 299284 101773
rect 299318 101745 299346 101773
rect 299380 101745 299408 101773
rect 299442 101745 299470 101773
rect 299256 92931 299284 92959
rect 299318 92931 299346 92959
rect 299380 92931 299408 92959
rect 299442 92931 299470 92959
rect 299256 92869 299284 92897
rect 299318 92869 299346 92897
rect 299380 92869 299408 92897
rect 299442 92869 299470 92897
rect 299256 92807 299284 92835
rect 299318 92807 299346 92835
rect 299380 92807 299408 92835
rect 299442 92807 299470 92835
rect 299256 92745 299284 92773
rect 299318 92745 299346 92773
rect 299380 92745 299408 92773
rect 299442 92745 299470 92773
rect 299256 83931 299284 83959
rect 299318 83931 299346 83959
rect 299380 83931 299408 83959
rect 299442 83931 299470 83959
rect 299256 83869 299284 83897
rect 299318 83869 299346 83897
rect 299380 83869 299408 83897
rect 299442 83869 299470 83897
rect 299256 83807 299284 83835
rect 299318 83807 299346 83835
rect 299380 83807 299408 83835
rect 299442 83807 299470 83835
rect 299256 83745 299284 83773
rect 299318 83745 299346 83773
rect 299380 83745 299408 83773
rect 299442 83745 299470 83773
rect 299256 74931 299284 74959
rect 299318 74931 299346 74959
rect 299380 74931 299408 74959
rect 299442 74931 299470 74959
rect 299256 74869 299284 74897
rect 299318 74869 299346 74897
rect 299380 74869 299408 74897
rect 299442 74869 299470 74897
rect 299256 74807 299284 74835
rect 299318 74807 299346 74835
rect 299380 74807 299408 74835
rect 299442 74807 299470 74835
rect 299256 74745 299284 74773
rect 299318 74745 299346 74773
rect 299380 74745 299408 74773
rect 299442 74745 299470 74773
rect 299256 65931 299284 65959
rect 299318 65931 299346 65959
rect 299380 65931 299408 65959
rect 299442 65931 299470 65959
rect 299256 65869 299284 65897
rect 299318 65869 299346 65897
rect 299380 65869 299408 65897
rect 299442 65869 299470 65897
rect 299256 65807 299284 65835
rect 299318 65807 299346 65835
rect 299380 65807 299408 65835
rect 299442 65807 299470 65835
rect 299256 65745 299284 65773
rect 299318 65745 299346 65773
rect 299380 65745 299408 65773
rect 299442 65745 299470 65773
rect 299256 56931 299284 56959
rect 299318 56931 299346 56959
rect 299380 56931 299408 56959
rect 299442 56931 299470 56959
rect 299256 56869 299284 56897
rect 299318 56869 299346 56897
rect 299380 56869 299408 56897
rect 299442 56869 299470 56897
rect 299256 56807 299284 56835
rect 299318 56807 299346 56835
rect 299380 56807 299408 56835
rect 299442 56807 299470 56835
rect 299256 56745 299284 56773
rect 299318 56745 299346 56773
rect 299380 56745 299408 56773
rect 299442 56745 299470 56773
rect 299256 47931 299284 47959
rect 299318 47931 299346 47959
rect 299380 47931 299408 47959
rect 299442 47931 299470 47959
rect 299256 47869 299284 47897
rect 299318 47869 299346 47897
rect 299380 47869 299408 47897
rect 299442 47869 299470 47897
rect 299256 47807 299284 47835
rect 299318 47807 299346 47835
rect 299380 47807 299408 47835
rect 299442 47807 299470 47835
rect 299256 47745 299284 47773
rect 299318 47745 299346 47773
rect 299380 47745 299408 47773
rect 299442 47745 299470 47773
rect 299256 38931 299284 38959
rect 299318 38931 299346 38959
rect 299380 38931 299408 38959
rect 299442 38931 299470 38959
rect 299256 38869 299284 38897
rect 299318 38869 299346 38897
rect 299380 38869 299408 38897
rect 299442 38869 299470 38897
rect 299256 38807 299284 38835
rect 299318 38807 299346 38835
rect 299380 38807 299408 38835
rect 299442 38807 299470 38835
rect 299256 38745 299284 38773
rect 299318 38745 299346 38773
rect 299380 38745 299408 38773
rect 299442 38745 299470 38773
rect 299256 29931 299284 29959
rect 299318 29931 299346 29959
rect 299380 29931 299408 29959
rect 299442 29931 299470 29959
rect 299256 29869 299284 29897
rect 299318 29869 299346 29897
rect 299380 29869 299408 29897
rect 299442 29869 299470 29897
rect 299256 29807 299284 29835
rect 299318 29807 299346 29835
rect 299380 29807 299408 29835
rect 299442 29807 299470 29835
rect 299256 29745 299284 29773
rect 299318 29745 299346 29773
rect 299380 29745 299408 29773
rect 299442 29745 299470 29773
rect 299256 20931 299284 20959
rect 299318 20931 299346 20959
rect 299380 20931 299408 20959
rect 299442 20931 299470 20959
rect 299256 20869 299284 20897
rect 299318 20869 299346 20897
rect 299380 20869 299408 20897
rect 299442 20869 299470 20897
rect 299256 20807 299284 20835
rect 299318 20807 299346 20835
rect 299380 20807 299408 20835
rect 299442 20807 299470 20835
rect 299256 20745 299284 20773
rect 299318 20745 299346 20773
rect 299380 20745 299408 20773
rect 299442 20745 299470 20773
rect 299256 11931 299284 11959
rect 299318 11931 299346 11959
rect 299380 11931 299408 11959
rect 299442 11931 299470 11959
rect 299256 11869 299284 11897
rect 299318 11869 299346 11897
rect 299380 11869 299408 11897
rect 299442 11869 299470 11897
rect 299256 11807 299284 11835
rect 299318 11807 299346 11835
rect 299380 11807 299408 11835
rect 299442 11807 299470 11835
rect 299256 11745 299284 11773
rect 299318 11745 299346 11773
rect 299380 11745 299408 11773
rect 299442 11745 299470 11773
rect 299256 2931 299284 2959
rect 299318 2931 299346 2959
rect 299380 2931 299408 2959
rect 299442 2931 299470 2959
rect 299256 2869 299284 2897
rect 299318 2869 299346 2897
rect 299380 2869 299408 2897
rect 299442 2869 299470 2897
rect 299256 2807 299284 2835
rect 299318 2807 299346 2835
rect 299380 2807 299408 2835
rect 299442 2807 299470 2835
rect 299256 2745 299284 2773
rect 299318 2745 299346 2773
rect 299380 2745 299408 2773
rect 299442 2745 299470 2773
rect 299256 876 299284 904
rect 299318 876 299346 904
rect 299380 876 299408 904
rect 299442 876 299470 904
rect 299256 814 299284 842
rect 299318 814 299346 842
rect 299380 814 299408 842
rect 299442 814 299470 842
rect 299256 752 299284 780
rect 299318 752 299346 780
rect 299380 752 299408 780
rect 299442 752 299470 780
rect 299256 690 299284 718
rect 299318 690 299346 718
rect 299380 690 299408 718
rect 299442 690 299470 718
rect 299736 293931 299764 293959
rect 299798 293931 299826 293959
rect 299860 293931 299888 293959
rect 299922 293931 299950 293959
rect 299736 293869 299764 293897
rect 299798 293869 299826 293897
rect 299860 293869 299888 293897
rect 299922 293869 299950 293897
rect 299736 293807 299764 293835
rect 299798 293807 299826 293835
rect 299860 293807 299888 293835
rect 299922 293807 299950 293835
rect 299736 293745 299764 293773
rect 299798 293745 299826 293773
rect 299860 293745 299888 293773
rect 299922 293745 299950 293773
rect 299736 284931 299764 284959
rect 299798 284931 299826 284959
rect 299860 284931 299888 284959
rect 299922 284931 299950 284959
rect 299736 284869 299764 284897
rect 299798 284869 299826 284897
rect 299860 284869 299888 284897
rect 299922 284869 299950 284897
rect 299736 284807 299764 284835
rect 299798 284807 299826 284835
rect 299860 284807 299888 284835
rect 299922 284807 299950 284835
rect 299736 284745 299764 284773
rect 299798 284745 299826 284773
rect 299860 284745 299888 284773
rect 299922 284745 299950 284773
rect 299736 275931 299764 275959
rect 299798 275931 299826 275959
rect 299860 275931 299888 275959
rect 299922 275931 299950 275959
rect 299736 275869 299764 275897
rect 299798 275869 299826 275897
rect 299860 275869 299888 275897
rect 299922 275869 299950 275897
rect 299736 275807 299764 275835
rect 299798 275807 299826 275835
rect 299860 275807 299888 275835
rect 299922 275807 299950 275835
rect 299736 275745 299764 275773
rect 299798 275745 299826 275773
rect 299860 275745 299888 275773
rect 299922 275745 299950 275773
rect 299736 266931 299764 266959
rect 299798 266931 299826 266959
rect 299860 266931 299888 266959
rect 299922 266931 299950 266959
rect 299736 266869 299764 266897
rect 299798 266869 299826 266897
rect 299860 266869 299888 266897
rect 299922 266869 299950 266897
rect 299736 266807 299764 266835
rect 299798 266807 299826 266835
rect 299860 266807 299888 266835
rect 299922 266807 299950 266835
rect 299736 266745 299764 266773
rect 299798 266745 299826 266773
rect 299860 266745 299888 266773
rect 299922 266745 299950 266773
rect 299736 257931 299764 257959
rect 299798 257931 299826 257959
rect 299860 257931 299888 257959
rect 299922 257931 299950 257959
rect 299736 257869 299764 257897
rect 299798 257869 299826 257897
rect 299860 257869 299888 257897
rect 299922 257869 299950 257897
rect 299736 257807 299764 257835
rect 299798 257807 299826 257835
rect 299860 257807 299888 257835
rect 299922 257807 299950 257835
rect 299736 257745 299764 257773
rect 299798 257745 299826 257773
rect 299860 257745 299888 257773
rect 299922 257745 299950 257773
rect 299736 248931 299764 248959
rect 299798 248931 299826 248959
rect 299860 248931 299888 248959
rect 299922 248931 299950 248959
rect 299736 248869 299764 248897
rect 299798 248869 299826 248897
rect 299860 248869 299888 248897
rect 299922 248869 299950 248897
rect 299736 248807 299764 248835
rect 299798 248807 299826 248835
rect 299860 248807 299888 248835
rect 299922 248807 299950 248835
rect 299736 248745 299764 248773
rect 299798 248745 299826 248773
rect 299860 248745 299888 248773
rect 299922 248745 299950 248773
rect 299736 239931 299764 239959
rect 299798 239931 299826 239959
rect 299860 239931 299888 239959
rect 299922 239931 299950 239959
rect 299736 239869 299764 239897
rect 299798 239869 299826 239897
rect 299860 239869 299888 239897
rect 299922 239869 299950 239897
rect 299736 239807 299764 239835
rect 299798 239807 299826 239835
rect 299860 239807 299888 239835
rect 299922 239807 299950 239835
rect 299736 239745 299764 239773
rect 299798 239745 299826 239773
rect 299860 239745 299888 239773
rect 299922 239745 299950 239773
rect 299736 230931 299764 230959
rect 299798 230931 299826 230959
rect 299860 230931 299888 230959
rect 299922 230931 299950 230959
rect 299736 230869 299764 230897
rect 299798 230869 299826 230897
rect 299860 230869 299888 230897
rect 299922 230869 299950 230897
rect 299736 230807 299764 230835
rect 299798 230807 299826 230835
rect 299860 230807 299888 230835
rect 299922 230807 299950 230835
rect 299736 230745 299764 230773
rect 299798 230745 299826 230773
rect 299860 230745 299888 230773
rect 299922 230745 299950 230773
rect 299736 221931 299764 221959
rect 299798 221931 299826 221959
rect 299860 221931 299888 221959
rect 299922 221931 299950 221959
rect 299736 221869 299764 221897
rect 299798 221869 299826 221897
rect 299860 221869 299888 221897
rect 299922 221869 299950 221897
rect 299736 221807 299764 221835
rect 299798 221807 299826 221835
rect 299860 221807 299888 221835
rect 299922 221807 299950 221835
rect 299736 221745 299764 221773
rect 299798 221745 299826 221773
rect 299860 221745 299888 221773
rect 299922 221745 299950 221773
rect 299736 212931 299764 212959
rect 299798 212931 299826 212959
rect 299860 212931 299888 212959
rect 299922 212931 299950 212959
rect 299736 212869 299764 212897
rect 299798 212869 299826 212897
rect 299860 212869 299888 212897
rect 299922 212869 299950 212897
rect 299736 212807 299764 212835
rect 299798 212807 299826 212835
rect 299860 212807 299888 212835
rect 299922 212807 299950 212835
rect 299736 212745 299764 212773
rect 299798 212745 299826 212773
rect 299860 212745 299888 212773
rect 299922 212745 299950 212773
rect 299736 203931 299764 203959
rect 299798 203931 299826 203959
rect 299860 203931 299888 203959
rect 299922 203931 299950 203959
rect 299736 203869 299764 203897
rect 299798 203869 299826 203897
rect 299860 203869 299888 203897
rect 299922 203869 299950 203897
rect 299736 203807 299764 203835
rect 299798 203807 299826 203835
rect 299860 203807 299888 203835
rect 299922 203807 299950 203835
rect 299736 203745 299764 203773
rect 299798 203745 299826 203773
rect 299860 203745 299888 203773
rect 299922 203745 299950 203773
rect 299736 194931 299764 194959
rect 299798 194931 299826 194959
rect 299860 194931 299888 194959
rect 299922 194931 299950 194959
rect 299736 194869 299764 194897
rect 299798 194869 299826 194897
rect 299860 194869 299888 194897
rect 299922 194869 299950 194897
rect 299736 194807 299764 194835
rect 299798 194807 299826 194835
rect 299860 194807 299888 194835
rect 299922 194807 299950 194835
rect 299736 194745 299764 194773
rect 299798 194745 299826 194773
rect 299860 194745 299888 194773
rect 299922 194745 299950 194773
rect 299736 185931 299764 185959
rect 299798 185931 299826 185959
rect 299860 185931 299888 185959
rect 299922 185931 299950 185959
rect 299736 185869 299764 185897
rect 299798 185869 299826 185897
rect 299860 185869 299888 185897
rect 299922 185869 299950 185897
rect 299736 185807 299764 185835
rect 299798 185807 299826 185835
rect 299860 185807 299888 185835
rect 299922 185807 299950 185835
rect 299736 185745 299764 185773
rect 299798 185745 299826 185773
rect 299860 185745 299888 185773
rect 299922 185745 299950 185773
rect 299736 176931 299764 176959
rect 299798 176931 299826 176959
rect 299860 176931 299888 176959
rect 299922 176931 299950 176959
rect 299736 176869 299764 176897
rect 299798 176869 299826 176897
rect 299860 176869 299888 176897
rect 299922 176869 299950 176897
rect 299736 176807 299764 176835
rect 299798 176807 299826 176835
rect 299860 176807 299888 176835
rect 299922 176807 299950 176835
rect 299736 176745 299764 176773
rect 299798 176745 299826 176773
rect 299860 176745 299888 176773
rect 299922 176745 299950 176773
rect 299736 167931 299764 167959
rect 299798 167931 299826 167959
rect 299860 167931 299888 167959
rect 299922 167931 299950 167959
rect 299736 167869 299764 167897
rect 299798 167869 299826 167897
rect 299860 167869 299888 167897
rect 299922 167869 299950 167897
rect 299736 167807 299764 167835
rect 299798 167807 299826 167835
rect 299860 167807 299888 167835
rect 299922 167807 299950 167835
rect 299736 167745 299764 167773
rect 299798 167745 299826 167773
rect 299860 167745 299888 167773
rect 299922 167745 299950 167773
rect 299736 158931 299764 158959
rect 299798 158931 299826 158959
rect 299860 158931 299888 158959
rect 299922 158931 299950 158959
rect 299736 158869 299764 158897
rect 299798 158869 299826 158897
rect 299860 158869 299888 158897
rect 299922 158869 299950 158897
rect 299736 158807 299764 158835
rect 299798 158807 299826 158835
rect 299860 158807 299888 158835
rect 299922 158807 299950 158835
rect 299736 158745 299764 158773
rect 299798 158745 299826 158773
rect 299860 158745 299888 158773
rect 299922 158745 299950 158773
rect 299736 149931 299764 149959
rect 299798 149931 299826 149959
rect 299860 149931 299888 149959
rect 299922 149931 299950 149959
rect 299736 149869 299764 149897
rect 299798 149869 299826 149897
rect 299860 149869 299888 149897
rect 299922 149869 299950 149897
rect 299736 149807 299764 149835
rect 299798 149807 299826 149835
rect 299860 149807 299888 149835
rect 299922 149807 299950 149835
rect 299736 149745 299764 149773
rect 299798 149745 299826 149773
rect 299860 149745 299888 149773
rect 299922 149745 299950 149773
rect 299736 140931 299764 140959
rect 299798 140931 299826 140959
rect 299860 140931 299888 140959
rect 299922 140931 299950 140959
rect 299736 140869 299764 140897
rect 299798 140869 299826 140897
rect 299860 140869 299888 140897
rect 299922 140869 299950 140897
rect 299736 140807 299764 140835
rect 299798 140807 299826 140835
rect 299860 140807 299888 140835
rect 299922 140807 299950 140835
rect 299736 140745 299764 140773
rect 299798 140745 299826 140773
rect 299860 140745 299888 140773
rect 299922 140745 299950 140773
rect 299736 131931 299764 131959
rect 299798 131931 299826 131959
rect 299860 131931 299888 131959
rect 299922 131931 299950 131959
rect 299736 131869 299764 131897
rect 299798 131869 299826 131897
rect 299860 131869 299888 131897
rect 299922 131869 299950 131897
rect 299736 131807 299764 131835
rect 299798 131807 299826 131835
rect 299860 131807 299888 131835
rect 299922 131807 299950 131835
rect 299736 131745 299764 131773
rect 299798 131745 299826 131773
rect 299860 131745 299888 131773
rect 299922 131745 299950 131773
rect 299736 122931 299764 122959
rect 299798 122931 299826 122959
rect 299860 122931 299888 122959
rect 299922 122931 299950 122959
rect 299736 122869 299764 122897
rect 299798 122869 299826 122897
rect 299860 122869 299888 122897
rect 299922 122869 299950 122897
rect 299736 122807 299764 122835
rect 299798 122807 299826 122835
rect 299860 122807 299888 122835
rect 299922 122807 299950 122835
rect 299736 122745 299764 122773
rect 299798 122745 299826 122773
rect 299860 122745 299888 122773
rect 299922 122745 299950 122773
rect 299736 113931 299764 113959
rect 299798 113931 299826 113959
rect 299860 113931 299888 113959
rect 299922 113931 299950 113959
rect 299736 113869 299764 113897
rect 299798 113869 299826 113897
rect 299860 113869 299888 113897
rect 299922 113869 299950 113897
rect 299736 113807 299764 113835
rect 299798 113807 299826 113835
rect 299860 113807 299888 113835
rect 299922 113807 299950 113835
rect 299736 113745 299764 113773
rect 299798 113745 299826 113773
rect 299860 113745 299888 113773
rect 299922 113745 299950 113773
rect 299736 104931 299764 104959
rect 299798 104931 299826 104959
rect 299860 104931 299888 104959
rect 299922 104931 299950 104959
rect 299736 104869 299764 104897
rect 299798 104869 299826 104897
rect 299860 104869 299888 104897
rect 299922 104869 299950 104897
rect 299736 104807 299764 104835
rect 299798 104807 299826 104835
rect 299860 104807 299888 104835
rect 299922 104807 299950 104835
rect 299736 104745 299764 104773
rect 299798 104745 299826 104773
rect 299860 104745 299888 104773
rect 299922 104745 299950 104773
rect 299736 95931 299764 95959
rect 299798 95931 299826 95959
rect 299860 95931 299888 95959
rect 299922 95931 299950 95959
rect 299736 95869 299764 95897
rect 299798 95869 299826 95897
rect 299860 95869 299888 95897
rect 299922 95869 299950 95897
rect 299736 95807 299764 95835
rect 299798 95807 299826 95835
rect 299860 95807 299888 95835
rect 299922 95807 299950 95835
rect 299736 95745 299764 95773
rect 299798 95745 299826 95773
rect 299860 95745 299888 95773
rect 299922 95745 299950 95773
rect 299736 86931 299764 86959
rect 299798 86931 299826 86959
rect 299860 86931 299888 86959
rect 299922 86931 299950 86959
rect 299736 86869 299764 86897
rect 299798 86869 299826 86897
rect 299860 86869 299888 86897
rect 299922 86869 299950 86897
rect 299736 86807 299764 86835
rect 299798 86807 299826 86835
rect 299860 86807 299888 86835
rect 299922 86807 299950 86835
rect 299736 86745 299764 86773
rect 299798 86745 299826 86773
rect 299860 86745 299888 86773
rect 299922 86745 299950 86773
rect 299736 77931 299764 77959
rect 299798 77931 299826 77959
rect 299860 77931 299888 77959
rect 299922 77931 299950 77959
rect 299736 77869 299764 77897
rect 299798 77869 299826 77897
rect 299860 77869 299888 77897
rect 299922 77869 299950 77897
rect 299736 77807 299764 77835
rect 299798 77807 299826 77835
rect 299860 77807 299888 77835
rect 299922 77807 299950 77835
rect 299736 77745 299764 77773
rect 299798 77745 299826 77773
rect 299860 77745 299888 77773
rect 299922 77745 299950 77773
rect 299736 68931 299764 68959
rect 299798 68931 299826 68959
rect 299860 68931 299888 68959
rect 299922 68931 299950 68959
rect 299736 68869 299764 68897
rect 299798 68869 299826 68897
rect 299860 68869 299888 68897
rect 299922 68869 299950 68897
rect 299736 68807 299764 68835
rect 299798 68807 299826 68835
rect 299860 68807 299888 68835
rect 299922 68807 299950 68835
rect 299736 68745 299764 68773
rect 299798 68745 299826 68773
rect 299860 68745 299888 68773
rect 299922 68745 299950 68773
rect 299736 59931 299764 59959
rect 299798 59931 299826 59959
rect 299860 59931 299888 59959
rect 299922 59931 299950 59959
rect 299736 59869 299764 59897
rect 299798 59869 299826 59897
rect 299860 59869 299888 59897
rect 299922 59869 299950 59897
rect 299736 59807 299764 59835
rect 299798 59807 299826 59835
rect 299860 59807 299888 59835
rect 299922 59807 299950 59835
rect 299736 59745 299764 59773
rect 299798 59745 299826 59773
rect 299860 59745 299888 59773
rect 299922 59745 299950 59773
rect 299736 50931 299764 50959
rect 299798 50931 299826 50959
rect 299860 50931 299888 50959
rect 299922 50931 299950 50959
rect 299736 50869 299764 50897
rect 299798 50869 299826 50897
rect 299860 50869 299888 50897
rect 299922 50869 299950 50897
rect 299736 50807 299764 50835
rect 299798 50807 299826 50835
rect 299860 50807 299888 50835
rect 299922 50807 299950 50835
rect 299736 50745 299764 50773
rect 299798 50745 299826 50773
rect 299860 50745 299888 50773
rect 299922 50745 299950 50773
rect 299736 41931 299764 41959
rect 299798 41931 299826 41959
rect 299860 41931 299888 41959
rect 299922 41931 299950 41959
rect 299736 41869 299764 41897
rect 299798 41869 299826 41897
rect 299860 41869 299888 41897
rect 299922 41869 299950 41897
rect 299736 41807 299764 41835
rect 299798 41807 299826 41835
rect 299860 41807 299888 41835
rect 299922 41807 299950 41835
rect 299736 41745 299764 41773
rect 299798 41745 299826 41773
rect 299860 41745 299888 41773
rect 299922 41745 299950 41773
rect 299736 32931 299764 32959
rect 299798 32931 299826 32959
rect 299860 32931 299888 32959
rect 299922 32931 299950 32959
rect 299736 32869 299764 32897
rect 299798 32869 299826 32897
rect 299860 32869 299888 32897
rect 299922 32869 299950 32897
rect 299736 32807 299764 32835
rect 299798 32807 299826 32835
rect 299860 32807 299888 32835
rect 299922 32807 299950 32835
rect 299736 32745 299764 32773
rect 299798 32745 299826 32773
rect 299860 32745 299888 32773
rect 299922 32745 299950 32773
rect 299736 23931 299764 23959
rect 299798 23931 299826 23959
rect 299860 23931 299888 23959
rect 299922 23931 299950 23959
rect 299736 23869 299764 23897
rect 299798 23869 299826 23897
rect 299860 23869 299888 23897
rect 299922 23869 299950 23897
rect 299736 23807 299764 23835
rect 299798 23807 299826 23835
rect 299860 23807 299888 23835
rect 299922 23807 299950 23835
rect 299736 23745 299764 23773
rect 299798 23745 299826 23773
rect 299860 23745 299888 23773
rect 299922 23745 299950 23773
rect 299736 14931 299764 14959
rect 299798 14931 299826 14959
rect 299860 14931 299888 14959
rect 299922 14931 299950 14959
rect 299736 14869 299764 14897
rect 299798 14869 299826 14897
rect 299860 14869 299888 14897
rect 299922 14869 299950 14897
rect 299736 14807 299764 14835
rect 299798 14807 299826 14835
rect 299860 14807 299888 14835
rect 299922 14807 299950 14835
rect 299736 14745 299764 14773
rect 299798 14745 299826 14773
rect 299860 14745 299888 14773
rect 299922 14745 299950 14773
rect 299736 5931 299764 5959
rect 299798 5931 299826 5959
rect 299860 5931 299888 5959
rect 299922 5931 299950 5959
rect 299736 5869 299764 5897
rect 299798 5869 299826 5897
rect 299860 5869 299888 5897
rect 299922 5869 299950 5897
rect 299736 5807 299764 5835
rect 299798 5807 299826 5835
rect 299860 5807 299888 5835
rect 299922 5807 299950 5835
rect 299736 5745 299764 5773
rect 299798 5745 299826 5773
rect 299860 5745 299888 5773
rect 299922 5745 299950 5773
rect 292437 396 292465 424
rect 292499 396 292527 424
rect 292561 396 292589 424
rect 292623 396 292651 424
rect 292437 334 292465 362
rect 292499 334 292527 362
rect 292561 334 292589 362
rect 292623 334 292651 362
rect 292437 272 292465 300
rect 292499 272 292527 300
rect 292561 272 292589 300
rect 292623 272 292651 300
rect 292437 210 292465 238
rect 292499 210 292527 238
rect 292561 210 292589 238
rect 292623 210 292651 238
rect 299736 396 299764 424
rect 299798 396 299826 424
rect 299860 396 299888 424
rect 299922 396 299950 424
rect 299736 334 299764 362
rect 299798 334 299826 362
rect 299860 334 299888 362
rect 299922 334 299950 362
rect 299736 272 299764 300
rect 299798 272 299826 300
rect 299860 272 299888 300
rect 299922 272 299950 300
rect 299736 210 299764 238
rect 299798 210 299826 238
rect 299860 210 299888 238
rect 299922 210 299950 238
<< metal5 >>
rect -6 299670 299998 299718
rect -6 299642 42 299670
rect 70 299642 104 299670
rect 132 299642 166 299670
rect 194 299642 228 299670
rect 256 299642 4437 299670
rect 4465 299642 4499 299670
rect 4527 299642 4561 299670
rect 4589 299642 4623 299670
rect 4651 299642 13437 299670
rect 13465 299642 13499 299670
rect 13527 299642 13561 299670
rect 13589 299642 13623 299670
rect 13651 299642 22437 299670
rect 22465 299642 22499 299670
rect 22527 299642 22561 299670
rect 22589 299642 22623 299670
rect 22651 299642 31437 299670
rect 31465 299642 31499 299670
rect 31527 299642 31561 299670
rect 31589 299642 31623 299670
rect 31651 299642 40437 299670
rect 40465 299642 40499 299670
rect 40527 299642 40561 299670
rect 40589 299642 40623 299670
rect 40651 299642 49437 299670
rect 49465 299642 49499 299670
rect 49527 299642 49561 299670
rect 49589 299642 49623 299670
rect 49651 299642 58437 299670
rect 58465 299642 58499 299670
rect 58527 299642 58561 299670
rect 58589 299642 58623 299670
rect 58651 299642 67437 299670
rect 67465 299642 67499 299670
rect 67527 299642 67561 299670
rect 67589 299642 67623 299670
rect 67651 299642 76437 299670
rect 76465 299642 76499 299670
rect 76527 299642 76561 299670
rect 76589 299642 76623 299670
rect 76651 299642 85437 299670
rect 85465 299642 85499 299670
rect 85527 299642 85561 299670
rect 85589 299642 85623 299670
rect 85651 299642 94437 299670
rect 94465 299642 94499 299670
rect 94527 299642 94561 299670
rect 94589 299642 94623 299670
rect 94651 299642 103437 299670
rect 103465 299642 103499 299670
rect 103527 299642 103561 299670
rect 103589 299642 103623 299670
rect 103651 299642 112437 299670
rect 112465 299642 112499 299670
rect 112527 299642 112561 299670
rect 112589 299642 112623 299670
rect 112651 299642 121437 299670
rect 121465 299642 121499 299670
rect 121527 299642 121561 299670
rect 121589 299642 121623 299670
rect 121651 299642 130437 299670
rect 130465 299642 130499 299670
rect 130527 299642 130561 299670
rect 130589 299642 130623 299670
rect 130651 299642 139437 299670
rect 139465 299642 139499 299670
rect 139527 299642 139561 299670
rect 139589 299642 139623 299670
rect 139651 299642 148437 299670
rect 148465 299642 148499 299670
rect 148527 299642 148561 299670
rect 148589 299642 148623 299670
rect 148651 299642 157437 299670
rect 157465 299642 157499 299670
rect 157527 299642 157561 299670
rect 157589 299642 157623 299670
rect 157651 299642 166437 299670
rect 166465 299642 166499 299670
rect 166527 299642 166561 299670
rect 166589 299642 166623 299670
rect 166651 299642 175437 299670
rect 175465 299642 175499 299670
rect 175527 299642 175561 299670
rect 175589 299642 175623 299670
rect 175651 299642 184437 299670
rect 184465 299642 184499 299670
rect 184527 299642 184561 299670
rect 184589 299642 184623 299670
rect 184651 299642 193437 299670
rect 193465 299642 193499 299670
rect 193527 299642 193561 299670
rect 193589 299642 193623 299670
rect 193651 299642 202437 299670
rect 202465 299642 202499 299670
rect 202527 299642 202561 299670
rect 202589 299642 202623 299670
rect 202651 299642 211437 299670
rect 211465 299642 211499 299670
rect 211527 299642 211561 299670
rect 211589 299642 211623 299670
rect 211651 299642 220437 299670
rect 220465 299642 220499 299670
rect 220527 299642 220561 299670
rect 220589 299642 220623 299670
rect 220651 299642 229437 299670
rect 229465 299642 229499 299670
rect 229527 299642 229561 299670
rect 229589 299642 229623 299670
rect 229651 299642 238437 299670
rect 238465 299642 238499 299670
rect 238527 299642 238561 299670
rect 238589 299642 238623 299670
rect 238651 299642 247437 299670
rect 247465 299642 247499 299670
rect 247527 299642 247561 299670
rect 247589 299642 247623 299670
rect 247651 299642 256437 299670
rect 256465 299642 256499 299670
rect 256527 299642 256561 299670
rect 256589 299642 256623 299670
rect 256651 299642 265437 299670
rect 265465 299642 265499 299670
rect 265527 299642 265561 299670
rect 265589 299642 265623 299670
rect 265651 299642 274437 299670
rect 274465 299642 274499 299670
rect 274527 299642 274561 299670
rect 274589 299642 274623 299670
rect 274651 299642 283437 299670
rect 283465 299642 283499 299670
rect 283527 299642 283561 299670
rect 283589 299642 283623 299670
rect 283651 299642 292437 299670
rect 292465 299642 292499 299670
rect 292527 299642 292561 299670
rect 292589 299642 292623 299670
rect 292651 299642 299736 299670
rect 299764 299642 299798 299670
rect 299826 299642 299860 299670
rect 299888 299642 299922 299670
rect 299950 299642 299998 299670
rect -6 299608 299998 299642
rect -6 299580 42 299608
rect 70 299580 104 299608
rect 132 299580 166 299608
rect 194 299580 228 299608
rect 256 299580 4437 299608
rect 4465 299580 4499 299608
rect 4527 299580 4561 299608
rect 4589 299580 4623 299608
rect 4651 299580 13437 299608
rect 13465 299580 13499 299608
rect 13527 299580 13561 299608
rect 13589 299580 13623 299608
rect 13651 299580 22437 299608
rect 22465 299580 22499 299608
rect 22527 299580 22561 299608
rect 22589 299580 22623 299608
rect 22651 299580 31437 299608
rect 31465 299580 31499 299608
rect 31527 299580 31561 299608
rect 31589 299580 31623 299608
rect 31651 299580 40437 299608
rect 40465 299580 40499 299608
rect 40527 299580 40561 299608
rect 40589 299580 40623 299608
rect 40651 299580 49437 299608
rect 49465 299580 49499 299608
rect 49527 299580 49561 299608
rect 49589 299580 49623 299608
rect 49651 299580 58437 299608
rect 58465 299580 58499 299608
rect 58527 299580 58561 299608
rect 58589 299580 58623 299608
rect 58651 299580 67437 299608
rect 67465 299580 67499 299608
rect 67527 299580 67561 299608
rect 67589 299580 67623 299608
rect 67651 299580 76437 299608
rect 76465 299580 76499 299608
rect 76527 299580 76561 299608
rect 76589 299580 76623 299608
rect 76651 299580 85437 299608
rect 85465 299580 85499 299608
rect 85527 299580 85561 299608
rect 85589 299580 85623 299608
rect 85651 299580 94437 299608
rect 94465 299580 94499 299608
rect 94527 299580 94561 299608
rect 94589 299580 94623 299608
rect 94651 299580 103437 299608
rect 103465 299580 103499 299608
rect 103527 299580 103561 299608
rect 103589 299580 103623 299608
rect 103651 299580 112437 299608
rect 112465 299580 112499 299608
rect 112527 299580 112561 299608
rect 112589 299580 112623 299608
rect 112651 299580 121437 299608
rect 121465 299580 121499 299608
rect 121527 299580 121561 299608
rect 121589 299580 121623 299608
rect 121651 299580 130437 299608
rect 130465 299580 130499 299608
rect 130527 299580 130561 299608
rect 130589 299580 130623 299608
rect 130651 299580 139437 299608
rect 139465 299580 139499 299608
rect 139527 299580 139561 299608
rect 139589 299580 139623 299608
rect 139651 299580 148437 299608
rect 148465 299580 148499 299608
rect 148527 299580 148561 299608
rect 148589 299580 148623 299608
rect 148651 299580 157437 299608
rect 157465 299580 157499 299608
rect 157527 299580 157561 299608
rect 157589 299580 157623 299608
rect 157651 299580 166437 299608
rect 166465 299580 166499 299608
rect 166527 299580 166561 299608
rect 166589 299580 166623 299608
rect 166651 299580 175437 299608
rect 175465 299580 175499 299608
rect 175527 299580 175561 299608
rect 175589 299580 175623 299608
rect 175651 299580 184437 299608
rect 184465 299580 184499 299608
rect 184527 299580 184561 299608
rect 184589 299580 184623 299608
rect 184651 299580 193437 299608
rect 193465 299580 193499 299608
rect 193527 299580 193561 299608
rect 193589 299580 193623 299608
rect 193651 299580 202437 299608
rect 202465 299580 202499 299608
rect 202527 299580 202561 299608
rect 202589 299580 202623 299608
rect 202651 299580 211437 299608
rect 211465 299580 211499 299608
rect 211527 299580 211561 299608
rect 211589 299580 211623 299608
rect 211651 299580 220437 299608
rect 220465 299580 220499 299608
rect 220527 299580 220561 299608
rect 220589 299580 220623 299608
rect 220651 299580 229437 299608
rect 229465 299580 229499 299608
rect 229527 299580 229561 299608
rect 229589 299580 229623 299608
rect 229651 299580 238437 299608
rect 238465 299580 238499 299608
rect 238527 299580 238561 299608
rect 238589 299580 238623 299608
rect 238651 299580 247437 299608
rect 247465 299580 247499 299608
rect 247527 299580 247561 299608
rect 247589 299580 247623 299608
rect 247651 299580 256437 299608
rect 256465 299580 256499 299608
rect 256527 299580 256561 299608
rect 256589 299580 256623 299608
rect 256651 299580 265437 299608
rect 265465 299580 265499 299608
rect 265527 299580 265561 299608
rect 265589 299580 265623 299608
rect 265651 299580 274437 299608
rect 274465 299580 274499 299608
rect 274527 299580 274561 299608
rect 274589 299580 274623 299608
rect 274651 299580 283437 299608
rect 283465 299580 283499 299608
rect 283527 299580 283561 299608
rect 283589 299580 283623 299608
rect 283651 299580 292437 299608
rect 292465 299580 292499 299608
rect 292527 299580 292561 299608
rect 292589 299580 292623 299608
rect 292651 299580 299736 299608
rect 299764 299580 299798 299608
rect 299826 299580 299860 299608
rect 299888 299580 299922 299608
rect 299950 299580 299998 299608
rect -6 299546 299998 299580
rect -6 299518 42 299546
rect 70 299518 104 299546
rect 132 299518 166 299546
rect 194 299518 228 299546
rect 256 299518 4437 299546
rect 4465 299518 4499 299546
rect 4527 299518 4561 299546
rect 4589 299518 4623 299546
rect 4651 299518 13437 299546
rect 13465 299518 13499 299546
rect 13527 299518 13561 299546
rect 13589 299518 13623 299546
rect 13651 299518 22437 299546
rect 22465 299518 22499 299546
rect 22527 299518 22561 299546
rect 22589 299518 22623 299546
rect 22651 299518 31437 299546
rect 31465 299518 31499 299546
rect 31527 299518 31561 299546
rect 31589 299518 31623 299546
rect 31651 299518 40437 299546
rect 40465 299518 40499 299546
rect 40527 299518 40561 299546
rect 40589 299518 40623 299546
rect 40651 299518 49437 299546
rect 49465 299518 49499 299546
rect 49527 299518 49561 299546
rect 49589 299518 49623 299546
rect 49651 299518 58437 299546
rect 58465 299518 58499 299546
rect 58527 299518 58561 299546
rect 58589 299518 58623 299546
rect 58651 299518 67437 299546
rect 67465 299518 67499 299546
rect 67527 299518 67561 299546
rect 67589 299518 67623 299546
rect 67651 299518 76437 299546
rect 76465 299518 76499 299546
rect 76527 299518 76561 299546
rect 76589 299518 76623 299546
rect 76651 299518 85437 299546
rect 85465 299518 85499 299546
rect 85527 299518 85561 299546
rect 85589 299518 85623 299546
rect 85651 299518 94437 299546
rect 94465 299518 94499 299546
rect 94527 299518 94561 299546
rect 94589 299518 94623 299546
rect 94651 299518 103437 299546
rect 103465 299518 103499 299546
rect 103527 299518 103561 299546
rect 103589 299518 103623 299546
rect 103651 299518 112437 299546
rect 112465 299518 112499 299546
rect 112527 299518 112561 299546
rect 112589 299518 112623 299546
rect 112651 299518 121437 299546
rect 121465 299518 121499 299546
rect 121527 299518 121561 299546
rect 121589 299518 121623 299546
rect 121651 299518 130437 299546
rect 130465 299518 130499 299546
rect 130527 299518 130561 299546
rect 130589 299518 130623 299546
rect 130651 299518 139437 299546
rect 139465 299518 139499 299546
rect 139527 299518 139561 299546
rect 139589 299518 139623 299546
rect 139651 299518 148437 299546
rect 148465 299518 148499 299546
rect 148527 299518 148561 299546
rect 148589 299518 148623 299546
rect 148651 299518 157437 299546
rect 157465 299518 157499 299546
rect 157527 299518 157561 299546
rect 157589 299518 157623 299546
rect 157651 299518 166437 299546
rect 166465 299518 166499 299546
rect 166527 299518 166561 299546
rect 166589 299518 166623 299546
rect 166651 299518 175437 299546
rect 175465 299518 175499 299546
rect 175527 299518 175561 299546
rect 175589 299518 175623 299546
rect 175651 299518 184437 299546
rect 184465 299518 184499 299546
rect 184527 299518 184561 299546
rect 184589 299518 184623 299546
rect 184651 299518 193437 299546
rect 193465 299518 193499 299546
rect 193527 299518 193561 299546
rect 193589 299518 193623 299546
rect 193651 299518 202437 299546
rect 202465 299518 202499 299546
rect 202527 299518 202561 299546
rect 202589 299518 202623 299546
rect 202651 299518 211437 299546
rect 211465 299518 211499 299546
rect 211527 299518 211561 299546
rect 211589 299518 211623 299546
rect 211651 299518 220437 299546
rect 220465 299518 220499 299546
rect 220527 299518 220561 299546
rect 220589 299518 220623 299546
rect 220651 299518 229437 299546
rect 229465 299518 229499 299546
rect 229527 299518 229561 299546
rect 229589 299518 229623 299546
rect 229651 299518 238437 299546
rect 238465 299518 238499 299546
rect 238527 299518 238561 299546
rect 238589 299518 238623 299546
rect 238651 299518 247437 299546
rect 247465 299518 247499 299546
rect 247527 299518 247561 299546
rect 247589 299518 247623 299546
rect 247651 299518 256437 299546
rect 256465 299518 256499 299546
rect 256527 299518 256561 299546
rect 256589 299518 256623 299546
rect 256651 299518 265437 299546
rect 265465 299518 265499 299546
rect 265527 299518 265561 299546
rect 265589 299518 265623 299546
rect 265651 299518 274437 299546
rect 274465 299518 274499 299546
rect 274527 299518 274561 299546
rect 274589 299518 274623 299546
rect 274651 299518 283437 299546
rect 283465 299518 283499 299546
rect 283527 299518 283561 299546
rect 283589 299518 283623 299546
rect 283651 299518 292437 299546
rect 292465 299518 292499 299546
rect 292527 299518 292561 299546
rect 292589 299518 292623 299546
rect 292651 299518 299736 299546
rect 299764 299518 299798 299546
rect 299826 299518 299860 299546
rect 299888 299518 299922 299546
rect 299950 299518 299998 299546
rect -6 299484 299998 299518
rect -6 299456 42 299484
rect 70 299456 104 299484
rect 132 299456 166 299484
rect 194 299456 228 299484
rect 256 299456 4437 299484
rect 4465 299456 4499 299484
rect 4527 299456 4561 299484
rect 4589 299456 4623 299484
rect 4651 299456 13437 299484
rect 13465 299456 13499 299484
rect 13527 299456 13561 299484
rect 13589 299456 13623 299484
rect 13651 299456 22437 299484
rect 22465 299456 22499 299484
rect 22527 299456 22561 299484
rect 22589 299456 22623 299484
rect 22651 299456 31437 299484
rect 31465 299456 31499 299484
rect 31527 299456 31561 299484
rect 31589 299456 31623 299484
rect 31651 299456 40437 299484
rect 40465 299456 40499 299484
rect 40527 299456 40561 299484
rect 40589 299456 40623 299484
rect 40651 299456 49437 299484
rect 49465 299456 49499 299484
rect 49527 299456 49561 299484
rect 49589 299456 49623 299484
rect 49651 299456 58437 299484
rect 58465 299456 58499 299484
rect 58527 299456 58561 299484
rect 58589 299456 58623 299484
rect 58651 299456 67437 299484
rect 67465 299456 67499 299484
rect 67527 299456 67561 299484
rect 67589 299456 67623 299484
rect 67651 299456 76437 299484
rect 76465 299456 76499 299484
rect 76527 299456 76561 299484
rect 76589 299456 76623 299484
rect 76651 299456 85437 299484
rect 85465 299456 85499 299484
rect 85527 299456 85561 299484
rect 85589 299456 85623 299484
rect 85651 299456 94437 299484
rect 94465 299456 94499 299484
rect 94527 299456 94561 299484
rect 94589 299456 94623 299484
rect 94651 299456 103437 299484
rect 103465 299456 103499 299484
rect 103527 299456 103561 299484
rect 103589 299456 103623 299484
rect 103651 299456 112437 299484
rect 112465 299456 112499 299484
rect 112527 299456 112561 299484
rect 112589 299456 112623 299484
rect 112651 299456 121437 299484
rect 121465 299456 121499 299484
rect 121527 299456 121561 299484
rect 121589 299456 121623 299484
rect 121651 299456 130437 299484
rect 130465 299456 130499 299484
rect 130527 299456 130561 299484
rect 130589 299456 130623 299484
rect 130651 299456 139437 299484
rect 139465 299456 139499 299484
rect 139527 299456 139561 299484
rect 139589 299456 139623 299484
rect 139651 299456 148437 299484
rect 148465 299456 148499 299484
rect 148527 299456 148561 299484
rect 148589 299456 148623 299484
rect 148651 299456 157437 299484
rect 157465 299456 157499 299484
rect 157527 299456 157561 299484
rect 157589 299456 157623 299484
rect 157651 299456 166437 299484
rect 166465 299456 166499 299484
rect 166527 299456 166561 299484
rect 166589 299456 166623 299484
rect 166651 299456 175437 299484
rect 175465 299456 175499 299484
rect 175527 299456 175561 299484
rect 175589 299456 175623 299484
rect 175651 299456 184437 299484
rect 184465 299456 184499 299484
rect 184527 299456 184561 299484
rect 184589 299456 184623 299484
rect 184651 299456 193437 299484
rect 193465 299456 193499 299484
rect 193527 299456 193561 299484
rect 193589 299456 193623 299484
rect 193651 299456 202437 299484
rect 202465 299456 202499 299484
rect 202527 299456 202561 299484
rect 202589 299456 202623 299484
rect 202651 299456 211437 299484
rect 211465 299456 211499 299484
rect 211527 299456 211561 299484
rect 211589 299456 211623 299484
rect 211651 299456 220437 299484
rect 220465 299456 220499 299484
rect 220527 299456 220561 299484
rect 220589 299456 220623 299484
rect 220651 299456 229437 299484
rect 229465 299456 229499 299484
rect 229527 299456 229561 299484
rect 229589 299456 229623 299484
rect 229651 299456 238437 299484
rect 238465 299456 238499 299484
rect 238527 299456 238561 299484
rect 238589 299456 238623 299484
rect 238651 299456 247437 299484
rect 247465 299456 247499 299484
rect 247527 299456 247561 299484
rect 247589 299456 247623 299484
rect 247651 299456 256437 299484
rect 256465 299456 256499 299484
rect 256527 299456 256561 299484
rect 256589 299456 256623 299484
rect 256651 299456 265437 299484
rect 265465 299456 265499 299484
rect 265527 299456 265561 299484
rect 265589 299456 265623 299484
rect 265651 299456 274437 299484
rect 274465 299456 274499 299484
rect 274527 299456 274561 299484
rect 274589 299456 274623 299484
rect 274651 299456 283437 299484
rect 283465 299456 283499 299484
rect 283527 299456 283561 299484
rect 283589 299456 283623 299484
rect 283651 299456 292437 299484
rect 292465 299456 292499 299484
rect 292527 299456 292561 299484
rect 292589 299456 292623 299484
rect 292651 299456 299736 299484
rect 299764 299456 299798 299484
rect 299826 299456 299860 299484
rect 299888 299456 299922 299484
rect 299950 299456 299998 299484
rect -6 299408 299998 299456
rect 474 299190 299518 299238
rect 474 299162 522 299190
rect 550 299162 584 299190
rect 612 299162 646 299190
rect 674 299162 708 299190
rect 736 299162 2577 299190
rect 2605 299162 2639 299190
rect 2667 299162 2701 299190
rect 2729 299162 2763 299190
rect 2791 299162 11577 299190
rect 11605 299162 11639 299190
rect 11667 299162 11701 299190
rect 11729 299162 11763 299190
rect 11791 299162 20577 299190
rect 20605 299162 20639 299190
rect 20667 299162 20701 299190
rect 20729 299162 20763 299190
rect 20791 299162 29577 299190
rect 29605 299162 29639 299190
rect 29667 299162 29701 299190
rect 29729 299162 29763 299190
rect 29791 299162 38577 299190
rect 38605 299162 38639 299190
rect 38667 299162 38701 299190
rect 38729 299162 38763 299190
rect 38791 299162 47577 299190
rect 47605 299162 47639 299190
rect 47667 299162 47701 299190
rect 47729 299162 47763 299190
rect 47791 299162 56577 299190
rect 56605 299162 56639 299190
rect 56667 299162 56701 299190
rect 56729 299162 56763 299190
rect 56791 299162 65577 299190
rect 65605 299162 65639 299190
rect 65667 299162 65701 299190
rect 65729 299162 65763 299190
rect 65791 299162 74577 299190
rect 74605 299162 74639 299190
rect 74667 299162 74701 299190
rect 74729 299162 74763 299190
rect 74791 299162 83577 299190
rect 83605 299162 83639 299190
rect 83667 299162 83701 299190
rect 83729 299162 83763 299190
rect 83791 299162 92577 299190
rect 92605 299162 92639 299190
rect 92667 299162 92701 299190
rect 92729 299162 92763 299190
rect 92791 299162 101577 299190
rect 101605 299162 101639 299190
rect 101667 299162 101701 299190
rect 101729 299162 101763 299190
rect 101791 299162 110577 299190
rect 110605 299162 110639 299190
rect 110667 299162 110701 299190
rect 110729 299162 110763 299190
rect 110791 299162 119577 299190
rect 119605 299162 119639 299190
rect 119667 299162 119701 299190
rect 119729 299162 119763 299190
rect 119791 299162 128577 299190
rect 128605 299162 128639 299190
rect 128667 299162 128701 299190
rect 128729 299162 128763 299190
rect 128791 299162 137577 299190
rect 137605 299162 137639 299190
rect 137667 299162 137701 299190
rect 137729 299162 137763 299190
rect 137791 299162 146577 299190
rect 146605 299162 146639 299190
rect 146667 299162 146701 299190
rect 146729 299162 146763 299190
rect 146791 299162 155577 299190
rect 155605 299162 155639 299190
rect 155667 299162 155701 299190
rect 155729 299162 155763 299190
rect 155791 299162 164577 299190
rect 164605 299162 164639 299190
rect 164667 299162 164701 299190
rect 164729 299162 164763 299190
rect 164791 299162 173577 299190
rect 173605 299162 173639 299190
rect 173667 299162 173701 299190
rect 173729 299162 173763 299190
rect 173791 299162 182577 299190
rect 182605 299162 182639 299190
rect 182667 299162 182701 299190
rect 182729 299162 182763 299190
rect 182791 299162 191577 299190
rect 191605 299162 191639 299190
rect 191667 299162 191701 299190
rect 191729 299162 191763 299190
rect 191791 299162 200577 299190
rect 200605 299162 200639 299190
rect 200667 299162 200701 299190
rect 200729 299162 200763 299190
rect 200791 299162 209577 299190
rect 209605 299162 209639 299190
rect 209667 299162 209701 299190
rect 209729 299162 209763 299190
rect 209791 299162 218577 299190
rect 218605 299162 218639 299190
rect 218667 299162 218701 299190
rect 218729 299162 218763 299190
rect 218791 299162 227577 299190
rect 227605 299162 227639 299190
rect 227667 299162 227701 299190
rect 227729 299162 227763 299190
rect 227791 299162 236577 299190
rect 236605 299162 236639 299190
rect 236667 299162 236701 299190
rect 236729 299162 236763 299190
rect 236791 299162 245577 299190
rect 245605 299162 245639 299190
rect 245667 299162 245701 299190
rect 245729 299162 245763 299190
rect 245791 299162 254577 299190
rect 254605 299162 254639 299190
rect 254667 299162 254701 299190
rect 254729 299162 254763 299190
rect 254791 299162 263577 299190
rect 263605 299162 263639 299190
rect 263667 299162 263701 299190
rect 263729 299162 263763 299190
rect 263791 299162 272577 299190
rect 272605 299162 272639 299190
rect 272667 299162 272701 299190
rect 272729 299162 272763 299190
rect 272791 299162 281577 299190
rect 281605 299162 281639 299190
rect 281667 299162 281701 299190
rect 281729 299162 281763 299190
rect 281791 299162 290577 299190
rect 290605 299162 290639 299190
rect 290667 299162 290701 299190
rect 290729 299162 290763 299190
rect 290791 299162 299256 299190
rect 299284 299162 299318 299190
rect 299346 299162 299380 299190
rect 299408 299162 299442 299190
rect 299470 299162 299518 299190
rect 474 299128 299518 299162
rect 474 299100 522 299128
rect 550 299100 584 299128
rect 612 299100 646 299128
rect 674 299100 708 299128
rect 736 299100 2577 299128
rect 2605 299100 2639 299128
rect 2667 299100 2701 299128
rect 2729 299100 2763 299128
rect 2791 299100 11577 299128
rect 11605 299100 11639 299128
rect 11667 299100 11701 299128
rect 11729 299100 11763 299128
rect 11791 299100 20577 299128
rect 20605 299100 20639 299128
rect 20667 299100 20701 299128
rect 20729 299100 20763 299128
rect 20791 299100 29577 299128
rect 29605 299100 29639 299128
rect 29667 299100 29701 299128
rect 29729 299100 29763 299128
rect 29791 299100 38577 299128
rect 38605 299100 38639 299128
rect 38667 299100 38701 299128
rect 38729 299100 38763 299128
rect 38791 299100 47577 299128
rect 47605 299100 47639 299128
rect 47667 299100 47701 299128
rect 47729 299100 47763 299128
rect 47791 299100 56577 299128
rect 56605 299100 56639 299128
rect 56667 299100 56701 299128
rect 56729 299100 56763 299128
rect 56791 299100 65577 299128
rect 65605 299100 65639 299128
rect 65667 299100 65701 299128
rect 65729 299100 65763 299128
rect 65791 299100 74577 299128
rect 74605 299100 74639 299128
rect 74667 299100 74701 299128
rect 74729 299100 74763 299128
rect 74791 299100 83577 299128
rect 83605 299100 83639 299128
rect 83667 299100 83701 299128
rect 83729 299100 83763 299128
rect 83791 299100 92577 299128
rect 92605 299100 92639 299128
rect 92667 299100 92701 299128
rect 92729 299100 92763 299128
rect 92791 299100 101577 299128
rect 101605 299100 101639 299128
rect 101667 299100 101701 299128
rect 101729 299100 101763 299128
rect 101791 299100 110577 299128
rect 110605 299100 110639 299128
rect 110667 299100 110701 299128
rect 110729 299100 110763 299128
rect 110791 299100 119577 299128
rect 119605 299100 119639 299128
rect 119667 299100 119701 299128
rect 119729 299100 119763 299128
rect 119791 299100 128577 299128
rect 128605 299100 128639 299128
rect 128667 299100 128701 299128
rect 128729 299100 128763 299128
rect 128791 299100 137577 299128
rect 137605 299100 137639 299128
rect 137667 299100 137701 299128
rect 137729 299100 137763 299128
rect 137791 299100 146577 299128
rect 146605 299100 146639 299128
rect 146667 299100 146701 299128
rect 146729 299100 146763 299128
rect 146791 299100 155577 299128
rect 155605 299100 155639 299128
rect 155667 299100 155701 299128
rect 155729 299100 155763 299128
rect 155791 299100 164577 299128
rect 164605 299100 164639 299128
rect 164667 299100 164701 299128
rect 164729 299100 164763 299128
rect 164791 299100 173577 299128
rect 173605 299100 173639 299128
rect 173667 299100 173701 299128
rect 173729 299100 173763 299128
rect 173791 299100 182577 299128
rect 182605 299100 182639 299128
rect 182667 299100 182701 299128
rect 182729 299100 182763 299128
rect 182791 299100 191577 299128
rect 191605 299100 191639 299128
rect 191667 299100 191701 299128
rect 191729 299100 191763 299128
rect 191791 299100 200577 299128
rect 200605 299100 200639 299128
rect 200667 299100 200701 299128
rect 200729 299100 200763 299128
rect 200791 299100 209577 299128
rect 209605 299100 209639 299128
rect 209667 299100 209701 299128
rect 209729 299100 209763 299128
rect 209791 299100 218577 299128
rect 218605 299100 218639 299128
rect 218667 299100 218701 299128
rect 218729 299100 218763 299128
rect 218791 299100 227577 299128
rect 227605 299100 227639 299128
rect 227667 299100 227701 299128
rect 227729 299100 227763 299128
rect 227791 299100 236577 299128
rect 236605 299100 236639 299128
rect 236667 299100 236701 299128
rect 236729 299100 236763 299128
rect 236791 299100 245577 299128
rect 245605 299100 245639 299128
rect 245667 299100 245701 299128
rect 245729 299100 245763 299128
rect 245791 299100 254577 299128
rect 254605 299100 254639 299128
rect 254667 299100 254701 299128
rect 254729 299100 254763 299128
rect 254791 299100 263577 299128
rect 263605 299100 263639 299128
rect 263667 299100 263701 299128
rect 263729 299100 263763 299128
rect 263791 299100 272577 299128
rect 272605 299100 272639 299128
rect 272667 299100 272701 299128
rect 272729 299100 272763 299128
rect 272791 299100 281577 299128
rect 281605 299100 281639 299128
rect 281667 299100 281701 299128
rect 281729 299100 281763 299128
rect 281791 299100 290577 299128
rect 290605 299100 290639 299128
rect 290667 299100 290701 299128
rect 290729 299100 290763 299128
rect 290791 299100 299256 299128
rect 299284 299100 299318 299128
rect 299346 299100 299380 299128
rect 299408 299100 299442 299128
rect 299470 299100 299518 299128
rect 474 299066 299518 299100
rect 474 299038 522 299066
rect 550 299038 584 299066
rect 612 299038 646 299066
rect 674 299038 708 299066
rect 736 299038 2577 299066
rect 2605 299038 2639 299066
rect 2667 299038 2701 299066
rect 2729 299038 2763 299066
rect 2791 299038 11577 299066
rect 11605 299038 11639 299066
rect 11667 299038 11701 299066
rect 11729 299038 11763 299066
rect 11791 299038 20577 299066
rect 20605 299038 20639 299066
rect 20667 299038 20701 299066
rect 20729 299038 20763 299066
rect 20791 299038 29577 299066
rect 29605 299038 29639 299066
rect 29667 299038 29701 299066
rect 29729 299038 29763 299066
rect 29791 299038 38577 299066
rect 38605 299038 38639 299066
rect 38667 299038 38701 299066
rect 38729 299038 38763 299066
rect 38791 299038 47577 299066
rect 47605 299038 47639 299066
rect 47667 299038 47701 299066
rect 47729 299038 47763 299066
rect 47791 299038 56577 299066
rect 56605 299038 56639 299066
rect 56667 299038 56701 299066
rect 56729 299038 56763 299066
rect 56791 299038 65577 299066
rect 65605 299038 65639 299066
rect 65667 299038 65701 299066
rect 65729 299038 65763 299066
rect 65791 299038 74577 299066
rect 74605 299038 74639 299066
rect 74667 299038 74701 299066
rect 74729 299038 74763 299066
rect 74791 299038 83577 299066
rect 83605 299038 83639 299066
rect 83667 299038 83701 299066
rect 83729 299038 83763 299066
rect 83791 299038 92577 299066
rect 92605 299038 92639 299066
rect 92667 299038 92701 299066
rect 92729 299038 92763 299066
rect 92791 299038 101577 299066
rect 101605 299038 101639 299066
rect 101667 299038 101701 299066
rect 101729 299038 101763 299066
rect 101791 299038 110577 299066
rect 110605 299038 110639 299066
rect 110667 299038 110701 299066
rect 110729 299038 110763 299066
rect 110791 299038 119577 299066
rect 119605 299038 119639 299066
rect 119667 299038 119701 299066
rect 119729 299038 119763 299066
rect 119791 299038 128577 299066
rect 128605 299038 128639 299066
rect 128667 299038 128701 299066
rect 128729 299038 128763 299066
rect 128791 299038 137577 299066
rect 137605 299038 137639 299066
rect 137667 299038 137701 299066
rect 137729 299038 137763 299066
rect 137791 299038 146577 299066
rect 146605 299038 146639 299066
rect 146667 299038 146701 299066
rect 146729 299038 146763 299066
rect 146791 299038 155577 299066
rect 155605 299038 155639 299066
rect 155667 299038 155701 299066
rect 155729 299038 155763 299066
rect 155791 299038 164577 299066
rect 164605 299038 164639 299066
rect 164667 299038 164701 299066
rect 164729 299038 164763 299066
rect 164791 299038 173577 299066
rect 173605 299038 173639 299066
rect 173667 299038 173701 299066
rect 173729 299038 173763 299066
rect 173791 299038 182577 299066
rect 182605 299038 182639 299066
rect 182667 299038 182701 299066
rect 182729 299038 182763 299066
rect 182791 299038 191577 299066
rect 191605 299038 191639 299066
rect 191667 299038 191701 299066
rect 191729 299038 191763 299066
rect 191791 299038 200577 299066
rect 200605 299038 200639 299066
rect 200667 299038 200701 299066
rect 200729 299038 200763 299066
rect 200791 299038 209577 299066
rect 209605 299038 209639 299066
rect 209667 299038 209701 299066
rect 209729 299038 209763 299066
rect 209791 299038 218577 299066
rect 218605 299038 218639 299066
rect 218667 299038 218701 299066
rect 218729 299038 218763 299066
rect 218791 299038 227577 299066
rect 227605 299038 227639 299066
rect 227667 299038 227701 299066
rect 227729 299038 227763 299066
rect 227791 299038 236577 299066
rect 236605 299038 236639 299066
rect 236667 299038 236701 299066
rect 236729 299038 236763 299066
rect 236791 299038 245577 299066
rect 245605 299038 245639 299066
rect 245667 299038 245701 299066
rect 245729 299038 245763 299066
rect 245791 299038 254577 299066
rect 254605 299038 254639 299066
rect 254667 299038 254701 299066
rect 254729 299038 254763 299066
rect 254791 299038 263577 299066
rect 263605 299038 263639 299066
rect 263667 299038 263701 299066
rect 263729 299038 263763 299066
rect 263791 299038 272577 299066
rect 272605 299038 272639 299066
rect 272667 299038 272701 299066
rect 272729 299038 272763 299066
rect 272791 299038 281577 299066
rect 281605 299038 281639 299066
rect 281667 299038 281701 299066
rect 281729 299038 281763 299066
rect 281791 299038 290577 299066
rect 290605 299038 290639 299066
rect 290667 299038 290701 299066
rect 290729 299038 290763 299066
rect 290791 299038 299256 299066
rect 299284 299038 299318 299066
rect 299346 299038 299380 299066
rect 299408 299038 299442 299066
rect 299470 299038 299518 299066
rect 474 299004 299518 299038
rect 474 298976 522 299004
rect 550 298976 584 299004
rect 612 298976 646 299004
rect 674 298976 708 299004
rect 736 298976 2577 299004
rect 2605 298976 2639 299004
rect 2667 298976 2701 299004
rect 2729 298976 2763 299004
rect 2791 298976 11577 299004
rect 11605 298976 11639 299004
rect 11667 298976 11701 299004
rect 11729 298976 11763 299004
rect 11791 298976 20577 299004
rect 20605 298976 20639 299004
rect 20667 298976 20701 299004
rect 20729 298976 20763 299004
rect 20791 298976 29577 299004
rect 29605 298976 29639 299004
rect 29667 298976 29701 299004
rect 29729 298976 29763 299004
rect 29791 298976 38577 299004
rect 38605 298976 38639 299004
rect 38667 298976 38701 299004
rect 38729 298976 38763 299004
rect 38791 298976 47577 299004
rect 47605 298976 47639 299004
rect 47667 298976 47701 299004
rect 47729 298976 47763 299004
rect 47791 298976 56577 299004
rect 56605 298976 56639 299004
rect 56667 298976 56701 299004
rect 56729 298976 56763 299004
rect 56791 298976 65577 299004
rect 65605 298976 65639 299004
rect 65667 298976 65701 299004
rect 65729 298976 65763 299004
rect 65791 298976 74577 299004
rect 74605 298976 74639 299004
rect 74667 298976 74701 299004
rect 74729 298976 74763 299004
rect 74791 298976 83577 299004
rect 83605 298976 83639 299004
rect 83667 298976 83701 299004
rect 83729 298976 83763 299004
rect 83791 298976 92577 299004
rect 92605 298976 92639 299004
rect 92667 298976 92701 299004
rect 92729 298976 92763 299004
rect 92791 298976 101577 299004
rect 101605 298976 101639 299004
rect 101667 298976 101701 299004
rect 101729 298976 101763 299004
rect 101791 298976 110577 299004
rect 110605 298976 110639 299004
rect 110667 298976 110701 299004
rect 110729 298976 110763 299004
rect 110791 298976 119577 299004
rect 119605 298976 119639 299004
rect 119667 298976 119701 299004
rect 119729 298976 119763 299004
rect 119791 298976 128577 299004
rect 128605 298976 128639 299004
rect 128667 298976 128701 299004
rect 128729 298976 128763 299004
rect 128791 298976 137577 299004
rect 137605 298976 137639 299004
rect 137667 298976 137701 299004
rect 137729 298976 137763 299004
rect 137791 298976 146577 299004
rect 146605 298976 146639 299004
rect 146667 298976 146701 299004
rect 146729 298976 146763 299004
rect 146791 298976 155577 299004
rect 155605 298976 155639 299004
rect 155667 298976 155701 299004
rect 155729 298976 155763 299004
rect 155791 298976 164577 299004
rect 164605 298976 164639 299004
rect 164667 298976 164701 299004
rect 164729 298976 164763 299004
rect 164791 298976 173577 299004
rect 173605 298976 173639 299004
rect 173667 298976 173701 299004
rect 173729 298976 173763 299004
rect 173791 298976 182577 299004
rect 182605 298976 182639 299004
rect 182667 298976 182701 299004
rect 182729 298976 182763 299004
rect 182791 298976 191577 299004
rect 191605 298976 191639 299004
rect 191667 298976 191701 299004
rect 191729 298976 191763 299004
rect 191791 298976 200577 299004
rect 200605 298976 200639 299004
rect 200667 298976 200701 299004
rect 200729 298976 200763 299004
rect 200791 298976 209577 299004
rect 209605 298976 209639 299004
rect 209667 298976 209701 299004
rect 209729 298976 209763 299004
rect 209791 298976 218577 299004
rect 218605 298976 218639 299004
rect 218667 298976 218701 299004
rect 218729 298976 218763 299004
rect 218791 298976 227577 299004
rect 227605 298976 227639 299004
rect 227667 298976 227701 299004
rect 227729 298976 227763 299004
rect 227791 298976 236577 299004
rect 236605 298976 236639 299004
rect 236667 298976 236701 299004
rect 236729 298976 236763 299004
rect 236791 298976 245577 299004
rect 245605 298976 245639 299004
rect 245667 298976 245701 299004
rect 245729 298976 245763 299004
rect 245791 298976 254577 299004
rect 254605 298976 254639 299004
rect 254667 298976 254701 299004
rect 254729 298976 254763 299004
rect 254791 298976 263577 299004
rect 263605 298976 263639 299004
rect 263667 298976 263701 299004
rect 263729 298976 263763 299004
rect 263791 298976 272577 299004
rect 272605 298976 272639 299004
rect 272667 298976 272701 299004
rect 272729 298976 272763 299004
rect 272791 298976 281577 299004
rect 281605 298976 281639 299004
rect 281667 298976 281701 299004
rect 281729 298976 281763 299004
rect 281791 298976 290577 299004
rect 290605 298976 290639 299004
rect 290667 298976 290701 299004
rect 290729 298976 290763 299004
rect 290791 298976 299256 299004
rect 299284 298976 299318 299004
rect 299346 298976 299380 299004
rect 299408 298976 299442 299004
rect 299470 298976 299518 299004
rect 474 298928 299518 298976
rect -6 293959 299998 294007
rect -6 293931 42 293959
rect 70 293931 104 293959
rect 132 293931 166 293959
rect 194 293931 228 293959
rect 256 293931 4437 293959
rect 4465 293931 4499 293959
rect 4527 293931 4561 293959
rect 4589 293931 4623 293959
rect 4651 293931 13437 293959
rect 13465 293931 13499 293959
rect 13527 293931 13561 293959
rect 13589 293931 13623 293959
rect 13651 293931 22437 293959
rect 22465 293931 22499 293959
rect 22527 293931 22561 293959
rect 22589 293931 22623 293959
rect 22651 293931 31437 293959
rect 31465 293931 31499 293959
rect 31527 293931 31561 293959
rect 31589 293931 31623 293959
rect 31651 293931 40437 293959
rect 40465 293931 40499 293959
rect 40527 293931 40561 293959
rect 40589 293931 40623 293959
rect 40651 293931 49437 293959
rect 49465 293931 49499 293959
rect 49527 293931 49561 293959
rect 49589 293931 49623 293959
rect 49651 293931 58437 293959
rect 58465 293931 58499 293959
rect 58527 293931 58561 293959
rect 58589 293931 58623 293959
rect 58651 293931 67437 293959
rect 67465 293931 67499 293959
rect 67527 293931 67561 293959
rect 67589 293931 67623 293959
rect 67651 293931 76437 293959
rect 76465 293931 76499 293959
rect 76527 293931 76561 293959
rect 76589 293931 76623 293959
rect 76651 293931 85437 293959
rect 85465 293931 85499 293959
rect 85527 293931 85561 293959
rect 85589 293931 85623 293959
rect 85651 293931 94437 293959
rect 94465 293931 94499 293959
rect 94527 293931 94561 293959
rect 94589 293931 94623 293959
rect 94651 293931 103437 293959
rect 103465 293931 103499 293959
rect 103527 293931 103561 293959
rect 103589 293931 103623 293959
rect 103651 293931 112437 293959
rect 112465 293931 112499 293959
rect 112527 293931 112561 293959
rect 112589 293931 112623 293959
rect 112651 293931 121437 293959
rect 121465 293931 121499 293959
rect 121527 293931 121561 293959
rect 121589 293931 121623 293959
rect 121651 293931 130437 293959
rect 130465 293931 130499 293959
rect 130527 293931 130561 293959
rect 130589 293931 130623 293959
rect 130651 293931 139437 293959
rect 139465 293931 139499 293959
rect 139527 293931 139561 293959
rect 139589 293931 139623 293959
rect 139651 293931 148437 293959
rect 148465 293931 148499 293959
rect 148527 293931 148561 293959
rect 148589 293931 148623 293959
rect 148651 293931 157437 293959
rect 157465 293931 157499 293959
rect 157527 293931 157561 293959
rect 157589 293931 157623 293959
rect 157651 293931 166437 293959
rect 166465 293931 166499 293959
rect 166527 293931 166561 293959
rect 166589 293931 166623 293959
rect 166651 293931 175437 293959
rect 175465 293931 175499 293959
rect 175527 293931 175561 293959
rect 175589 293931 175623 293959
rect 175651 293931 184437 293959
rect 184465 293931 184499 293959
rect 184527 293931 184561 293959
rect 184589 293931 184623 293959
rect 184651 293931 193437 293959
rect 193465 293931 193499 293959
rect 193527 293931 193561 293959
rect 193589 293931 193623 293959
rect 193651 293931 202437 293959
rect 202465 293931 202499 293959
rect 202527 293931 202561 293959
rect 202589 293931 202623 293959
rect 202651 293931 211437 293959
rect 211465 293931 211499 293959
rect 211527 293931 211561 293959
rect 211589 293931 211623 293959
rect 211651 293931 220437 293959
rect 220465 293931 220499 293959
rect 220527 293931 220561 293959
rect 220589 293931 220623 293959
rect 220651 293931 229437 293959
rect 229465 293931 229499 293959
rect 229527 293931 229561 293959
rect 229589 293931 229623 293959
rect 229651 293931 238437 293959
rect 238465 293931 238499 293959
rect 238527 293931 238561 293959
rect 238589 293931 238623 293959
rect 238651 293931 247437 293959
rect 247465 293931 247499 293959
rect 247527 293931 247561 293959
rect 247589 293931 247623 293959
rect 247651 293931 256437 293959
rect 256465 293931 256499 293959
rect 256527 293931 256561 293959
rect 256589 293931 256623 293959
rect 256651 293931 265437 293959
rect 265465 293931 265499 293959
rect 265527 293931 265561 293959
rect 265589 293931 265623 293959
rect 265651 293931 274437 293959
rect 274465 293931 274499 293959
rect 274527 293931 274561 293959
rect 274589 293931 274623 293959
rect 274651 293931 283437 293959
rect 283465 293931 283499 293959
rect 283527 293931 283561 293959
rect 283589 293931 283623 293959
rect 283651 293931 292437 293959
rect 292465 293931 292499 293959
rect 292527 293931 292561 293959
rect 292589 293931 292623 293959
rect 292651 293931 299736 293959
rect 299764 293931 299798 293959
rect 299826 293931 299860 293959
rect 299888 293931 299922 293959
rect 299950 293931 299998 293959
rect -6 293897 299998 293931
rect -6 293869 42 293897
rect 70 293869 104 293897
rect 132 293869 166 293897
rect 194 293869 228 293897
rect 256 293869 4437 293897
rect 4465 293869 4499 293897
rect 4527 293869 4561 293897
rect 4589 293869 4623 293897
rect 4651 293869 13437 293897
rect 13465 293869 13499 293897
rect 13527 293869 13561 293897
rect 13589 293869 13623 293897
rect 13651 293869 22437 293897
rect 22465 293869 22499 293897
rect 22527 293869 22561 293897
rect 22589 293869 22623 293897
rect 22651 293869 31437 293897
rect 31465 293869 31499 293897
rect 31527 293869 31561 293897
rect 31589 293869 31623 293897
rect 31651 293869 40437 293897
rect 40465 293869 40499 293897
rect 40527 293869 40561 293897
rect 40589 293869 40623 293897
rect 40651 293869 49437 293897
rect 49465 293869 49499 293897
rect 49527 293869 49561 293897
rect 49589 293869 49623 293897
rect 49651 293869 58437 293897
rect 58465 293869 58499 293897
rect 58527 293869 58561 293897
rect 58589 293869 58623 293897
rect 58651 293869 67437 293897
rect 67465 293869 67499 293897
rect 67527 293869 67561 293897
rect 67589 293869 67623 293897
rect 67651 293869 76437 293897
rect 76465 293869 76499 293897
rect 76527 293869 76561 293897
rect 76589 293869 76623 293897
rect 76651 293869 85437 293897
rect 85465 293869 85499 293897
rect 85527 293869 85561 293897
rect 85589 293869 85623 293897
rect 85651 293869 94437 293897
rect 94465 293869 94499 293897
rect 94527 293869 94561 293897
rect 94589 293869 94623 293897
rect 94651 293869 103437 293897
rect 103465 293869 103499 293897
rect 103527 293869 103561 293897
rect 103589 293869 103623 293897
rect 103651 293869 112437 293897
rect 112465 293869 112499 293897
rect 112527 293869 112561 293897
rect 112589 293869 112623 293897
rect 112651 293869 121437 293897
rect 121465 293869 121499 293897
rect 121527 293869 121561 293897
rect 121589 293869 121623 293897
rect 121651 293869 130437 293897
rect 130465 293869 130499 293897
rect 130527 293869 130561 293897
rect 130589 293869 130623 293897
rect 130651 293869 139437 293897
rect 139465 293869 139499 293897
rect 139527 293869 139561 293897
rect 139589 293869 139623 293897
rect 139651 293869 148437 293897
rect 148465 293869 148499 293897
rect 148527 293869 148561 293897
rect 148589 293869 148623 293897
rect 148651 293869 157437 293897
rect 157465 293869 157499 293897
rect 157527 293869 157561 293897
rect 157589 293869 157623 293897
rect 157651 293869 166437 293897
rect 166465 293869 166499 293897
rect 166527 293869 166561 293897
rect 166589 293869 166623 293897
rect 166651 293869 175437 293897
rect 175465 293869 175499 293897
rect 175527 293869 175561 293897
rect 175589 293869 175623 293897
rect 175651 293869 184437 293897
rect 184465 293869 184499 293897
rect 184527 293869 184561 293897
rect 184589 293869 184623 293897
rect 184651 293869 193437 293897
rect 193465 293869 193499 293897
rect 193527 293869 193561 293897
rect 193589 293869 193623 293897
rect 193651 293869 202437 293897
rect 202465 293869 202499 293897
rect 202527 293869 202561 293897
rect 202589 293869 202623 293897
rect 202651 293869 211437 293897
rect 211465 293869 211499 293897
rect 211527 293869 211561 293897
rect 211589 293869 211623 293897
rect 211651 293869 220437 293897
rect 220465 293869 220499 293897
rect 220527 293869 220561 293897
rect 220589 293869 220623 293897
rect 220651 293869 229437 293897
rect 229465 293869 229499 293897
rect 229527 293869 229561 293897
rect 229589 293869 229623 293897
rect 229651 293869 238437 293897
rect 238465 293869 238499 293897
rect 238527 293869 238561 293897
rect 238589 293869 238623 293897
rect 238651 293869 247437 293897
rect 247465 293869 247499 293897
rect 247527 293869 247561 293897
rect 247589 293869 247623 293897
rect 247651 293869 256437 293897
rect 256465 293869 256499 293897
rect 256527 293869 256561 293897
rect 256589 293869 256623 293897
rect 256651 293869 265437 293897
rect 265465 293869 265499 293897
rect 265527 293869 265561 293897
rect 265589 293869 265623 293897
rect 265651 293869 274437 293897
rect 274465 293869 274499 293897
rect 274527 293869 274561 293897
rect 274589 293869 274623 293897
rect 274651 293869 283437 293897
rect 283465 293869 283499 293897
rect 283527 293869 283561 293897
rect 283589 293869 283623 293897
rect 283651 293869 292437 293897
rect 292465 293869 292499 293897
rect 292527 293869 292561 293897
rect 292589 293869 292623 293897
rect 292651 293869 299736 293897
rect 299764 293869 299798 293897
rect 299826 293869 299860 293897
rect 299888 293869 299922 293897
rect 299950 293869 299998 293897
rect -6 293835 299998 293869
rect -6 293807 42 293835
rect 70 293807 104 293835
rect 132 293807 166 293835
rect 194 293807 228 293835
rect 256 293807 4437 293835
rect 4465 293807 4499 293835
rect 4527 293807 4561 293835
rect 4589 293807 4623 293835
rect 4651 293807 13437 293835
rect 13465 293807 13499 293835
rect 13527 293807 13561 293835
rect 13589 293807 13623 293835
rect 13651 293807 22437 293835
rect 22465 293807 22499 293835
rect 22527 293807 22561 293835
rect 22589 293807 22623 293835
rect 22651 293807 31437 293835
rect 31465 293807 31499 293835
rect 31527 293807 31561 293835
rect 31589 293807 31623 293835
rect 31651 293807 40437 293835
rect 40465 293807 40499 293835
rect 40527 293807 40561 293835
rect 40589 293807 40623 293835
rect 40651 293807 49437 293835
rect 49465 293807 49499 293835
rect 49527 293807 49561 293835
rect 49589 293807 49623 293835
rect 49651 293807 58437 293835
rect 58465 293807 58499 293835
rect 58527 293807 58561 293835
rect 58589 293807 58623 293835
rect 58651 293807 67437 293835
rect 67465 293807 67499 293835
rect 67527 293807 67561 293835
rect 67589 293807 67623 293835
rect 67651 293807 76437 293835
rect 76465 293807 76499 293835
rect 76527 293807 76561 293835
rect 76589 293807 76623 293835
rect 76651 293807 85437 293835
rect 85465 293807 85499 293835
rect 85527 293807 85561 293835
rect 85589 293807 85623 293835
rect 85651 293807 94437 293835
rect 94465 293807 94499 293835
rect 94527 293807 94561 293835
rect 94589 293807 94623 293835
rect 94651 293807 103437 293835
rect 103465 293807 103499 293835
rect 103527 293807 103561 293835
rect 103589 293807 103623 293835
rect 103651 293807 112437 293835
rect 112465 293807 112499 293835
rect 112527 293807 112561 293835
rect 112589 293807 112623 293835
rect 112651 293807 121437 293835
rect 121465 293807 121499 293835
rect 121527 293807 121561 293835
rect 121589 293807 121623 293835
rect 121651 293807 130437 293835
rect 130465 293807 130499 293835
rect 130527 293807 130561 293835
rect 130589 293807 130623 293835
rect 130651 293807 139437 293835
rect 139465 293807 139499 293835
rect 139527 293807 139561 293835
rect 139589 293807 139623 293835
rect 139651 293807 148437 293835
rect 148465 293807 148499 293835
rect 148527 293807 148561 293835
rect 148589 293807 148623 293835
rect 148651 293807 157437 293835
rect 157465 293807 157499 293835
rect 157527 293807 157561 293835
rect 157589 293807 157623 293835
rect 157651 293807 166437 293835
rect 166465 293807 166499 293835
rect 166527 293807 166561 293835
rect 166589 293807 166623 293835
rect 166651 293807 175437 293835
rect 175465 293807 175499 293835
rect 175527 293807 175561 293835
rect 175589 293807 175623 293835
rect 175651 293807 184437 293835
rect 184465 293807 184499 293835
rect 184527 293807 184561 293835
rect 184589 293807 184623 293835
rect 184651 293807 193437 293835
rect 193465 293807 193499 293835
rect 193527 293807 193561 293835
rect 193589 293807 193623 293835
rect 193651 293807 202437 293835
rect 202465 293807 202499 293835
rect 202527 293807 202561 293835
rect 202589 293807 202623 293835
rect 202651 293807 211437 293835
rect 211465 293807 211499 293835
rect 211527 293807 211561 293835
rect 211589 293807 211623 293835
rect 211651 293807 220437 293835
rect 220465 293807 220499 293835
rect 220527 293807 220561 293835
rect 220589 293807 220623 293835
rect 220651 293807 229437 293835
rect 229465 293807 229499 293835
rect 229527 293807 229561 293835
rect 229589 293807 229623 293835
rect 229651 293807 238437 293835
rect 238465 293807 238499 293835
rect 238527 293807 238561 293835
rect 238589 293807 238623 293835
rect 238651 293807 247437 293835
rect 247465 293807 247499 293835
rect 247527 293807 247561 293835
rect 247589 293807 247623 293835
rect 247651 293807 256437 293835
rect 256465 293807 256499 293835
rect 256527 293807 256561 293835
rect 256589 293807 256623 293835
rect 256651 293807 265437 293835
rect 265465 293807 265499 293835
rect 265527 293807 265561 293835
rect 265589 293807 265623 293835
rect 265651 293807 274437 293835
rect 274465 293807 274499 293835
rect 274527 293807 274561 293835
rect 274589 293807 274623 293835
rect 274651 293807 283437 293835
rect 283465 293807 283499 293835
rect 283527 293807 283561 293835
rect 283589 293807 283623 293835
rect 283651 293807 292437 293835
rect 292465 293807 292499 293835
rect 292527 293807 292561 293835
rect 292589 293807 292623 293835
rect 292651 293807 299736 293835
rect 299764 293807 299798 293835
rect 299826 293807 299860 293835
rect 299888 293807 299922 293835
rect 299950 293807 299998 293835
rect -6 293773 299998 293807
rect -6 293745 42 293773
rect 70 293745 104 293773
rect 132 293745 166 293773
rect 194 293745 228 293773
rect 256 293745 4437 293773
rect 4465 293745 4499 293773
rect 4527 293745 4561 293773
rect 4589 293745 4623 293773
rect 4651 293745 13437 293773
rect 13465 293745 13499 293773
rect 13527 293745 13561 293773
rect 13589 293745 13623 293773
rect 13651 293745 22437 293773
rect 22465 293745 22499 293773
rect 22527 293745 22561 293773
rect 22589 293745 22623 293773
rect 22651 293745 31437 293773
rect 31465 293745 31499 293773
rect 31527 293745 31561 293773
rect 31589 293745 31623 293773
rect 31651 293745 40437 293773
rect 40465 293745 40499 293773
rect 40527 293745 40561 293773
rect 40589 293745 40623 293773
rect 40651 293745 49437 293773
rect 49465 293745 49499 293773
rect 49527 293745 49561 293773
rect 49589 293745 49623 293773
rect 49651 293745 58437 293773
rect 58465 293745 58499 293773
rect 58527 293745 58561 293773
rect 58589 293745 58623 293773
rect 58651 293745 67437 293773
rect 67465 293745 67499 293773
rect 67527 293745 67561 293773
rect 67589 293745 67623 293773
rect 67651 293745 76437 293773
rect 76465 293745 76499 293773
rect 76527 293745 76561 293773
rect 76589 293745 76623 293773
rect 76651 293745 85437 293773
rect 85465 293745 85499 293773
rect 85527 293745 85561 293773
rect 85589 293745 85623 293773
rect 85651 293745 94437 293773
rect 94465 293745 94499 293773
rect 94527 293745 94561 293773
rect 94589 293745 94623 293773
rect 94651 293745 103437 293773
rect 103465 293745 103499 293773
rect 103527 293745 103561 293773
rect 103589 293745 103623 293773
rect 103651 293745 112437 293773
rect 112465 293745 112499 293773
rect 112527 293745 112561 293773
rect 112589 293745 112623 293773
rect 112651 293745 121437 293773
rect 121465 293745 121499 293773
rect 121527 293745 121561 293773
rect 121589 293745 121623 293773
rect 121651 293745 130437 293773
rect 130465 293745 130499 293773
rect 130527 293745 130561 293773
rect 130589 293745 130623 293773
rect 130651 293745 139437 293773
rect 139465 293745 139499 293773
rect 139527 293745 139561 293773
rect 139589 293745 139623 293773
rect 139651 293745 148437 293773
rect 148465 293745 148499 293773
rect 148527 293745 148561 293773
rect 148589 293745 148623 293773
rect 148651 293745 157437 293773
rect 157465 293745 157499 293773
rect 157527 293745 157561 293773
rect 157589 293745 157623 293773
rect 157651 293745 166437 293773
rect 166465 293745 166499 293773
rect 166527 293745 166561 293773
rect 166589 293745 166623 293773
rect 166651 293745 175437 293773
rect 175465 293745 175499 293773
rect 175527 293745 175561 293773
rect 175589 293745 175623 293773
rect 175651 293745 184437 293773
rect 184465 293745 184499 293773
rect 184527 293745 184561 293773
rect 184589 293745 184623 293773
rect 184651 293745 193437 293773
rect 193465 293745 193499 293773
rect 193527 293745 193561 293773
rect 193589 293745 193623 293773
rect 193651 293745 202437 293773
rect 202465 293745 202499 293773
rect 202527 293745 202561 293773
rect 202589 293745 202623 293773
rect 202651 293745 211437 293773
rect 211465 293745 211499 293773
rect 211527 293745 211561 293773
rect 211589 293745 211623 293773
rect 211651 293745 220437 293773
rect 220465 293745 220499 293773
rect 220527 293745 220561 293773
rect 220589 293745 220623 293773
rect 220651 293745 229437 293773
rect 229465 293745 229499 293773
rect 229527 293745 229561 293773
rect 229589 293745 229623 293773
rect 229651 293745 238437 293773
rect 238465 293745 238499 293773
rect 238527 293745 238561 293773
rect 238589 293745 238623 293773
rect 238651 293745 247437 293773
rect 247465 293745 247499 293773
rect 247527 293745 247561 293773
rect 247589 293745 247623 293773
rect 247651 293745 256437 293773
rect 256465 293745 256499 293773
rect 256527 293745 256561 293773
rect 256589 293745 256623 293773
rect 256651 293745 265437 293773
rect 265465 293745 265499 293773
rect 265527 293745 265561 293773
rect 265589 293745 265623 293773
rect 265651 293745 274437 293773
rect 274465 293745 274499 293773
rect 274527 293745 274561 293773
rect 274589 293745 274623 293773
rect 274651 293745 283437 293773
rect 283465 293745 283499 293773
rect 283527 293745 283561 293773
rect 283589 293745 283623 293773
rect 283651 293745 292437 293773
rect 292465 293745 292499 293773
rect 292527 293745 292561 293773
rect 292589 293745 292623 293773
rect 292651 293745 299736 293773
rect 299764 293745 299798 293773
rect 299826 293745 299860 293773
rect 299888 293745 299922 293773
rect 299950 293745 299998 293773
rect -6 293697 299998 293745
rect -6 290959 299998 291007
rect -6 290931 522 290959
rect 550 290931 584 290959
rect 612 290931 646 290959
rect 674 290931 708 290959
rect 736 290931 2577 290959
rect 2605 290931 2639 290959
rect 2667 290931 2701 290959
rect 2729 290931 2763 290959
rect 2791 290931 11577 290959
rect 11605 290931 11639 290959
rect 11667 290931 11701 290959
rect 11729 290931 11763 290959
rect 11791 290931 20577 290959
rect 20605 290931 20639 290959
rect 20667 290931 20701 290959
rect 20729 290931 20763 290959
rect 20791 290931 29577 290959
rect 29605 290931 29639 290959
rect 29667 290931 29701 290959
rect 29729 290931 29763 290959
rect 29791 290931 38577 290959
rect 38605 290931 38639 290959
rect 38667 290931 38701 290959
rect 38729 290931 38763 290959
rect 38791 290931 47577 290959
rect 47605 290931 47639 290959
rect 47667 290931 47701 290959
rect 47729 290931 47763 290959
rect 47791 290931 56577 290959
rect 56605 290931 56639 290959
rect 56667 290931 56701 290959
rect 56729 290931 56763 290959
rect 56791 290931 65577 290959
rect 65605 290931 65639 290959
rect 65667 290931 65701 290959
rect 65729 290931 65763 290959
rect 65791 290931 74577 290959
rect 74605 290931 74639 290959
rect 74667 290931 74701 290959
rect 74729 290931 74763 290959
rect 74791 290931 83577 290959
rect 83605 290931 83639 290959
rect 83667 290931 83701 290959
rect 83729 290931 83763 290959
rect 83791 290931 92577 290959
rect 92605 290931 92639 290959
rect 92667 290931 92701 290959
rect 92729 290931 92763 290959
rect 92791 290931 101577 290959
rect 101605 290931 101639 290959
rect 101667 290931 101701 290959
rect 101729 290931 101763 290959
rect 101791 290931 110577 290959
rect 110605 290931 110639 290959
rect 110667 290931 110701 290959
rect 110729 290931 110763 290959
rect 110791 290931 119577 290959
rect 119605 290931 119639 290959
rect 119667 290931 119701 290959
rect 119729 290931 119763 290959
rect 119791 290931 128577 290959
rect 128605 290931 128639 290959
rect 128667 290931 128701 290959
rect 128729 290931 128763 290959
rect 128791 290931 137577 290959
rect 137605 290931 137639 290959
rect 137667 290931 137701 290959
rect 137729 290931 137763 290959
rect 137791 290931 146577 290959
rect 146605 290931 146639 290959
rect 146667 290931 146701 290959
rect 146729 290931 146763 290959
rect 146791 290931 155577 290959
rect 155605 290931 155639 290959
rect 155667 290931 155701 290959
rect 155729 290931 155763 290959
rect 155791 290931 164577 290959
rect 164605 290931 164639 290959
rect 164667 290931 164701 290959
rect 164729 290931 164763 290959
rect 164791 290931 173577 290959
rect 173605 290931 173639 290959
rect 173667 290931 173701 290959
rect 173729 290931 173763 290959
rect 173791 290931 182577 290959
rect 182605 290931 182639 290959
rect 182667 290931 182701 290959
rect 182729 290931 182763 290959
rect 182791 290931 191577 290959
rect 191605 290931 191639 290959
rect 191667 290931 191701 290959
rect 191729 290931 191763 290959
rect 191791 290931 200577 290959
rect 200605 290931 200639 290959
rect 200667 290931 200701 290959
rect 200729 290931 200763 290959
rect 200791 290931 209577 290959
rect 209605 290931 209639 290959
rect 209667 290931 209701 290959
rect 209729 290931 209763 290959
rect 209791 290931 218577 290959
rect 218605 290931 218639 290959
rect 218667 290931 218701 290959
rect 218729 290931 218763 290959
rect 218791 290931 227577 290959
rect 227605 290931 227639 290959
rect 227667 290931 227701 290959
rect 227729 290931 227763 290959
rect 227791 290931 236577 290959
rect 236605 290931 236639 290959
rect 236667 290931 236701 290959
rect 236729 290931 236763 290959
rect 236791 290931 245577 290959
rect 245605 290931 245639 290959
rect 245667 290931 245701 290959
rect 245729 290931 245763 290959
rect 245791 290931 254577 290959
rect 254605 290931 254639 290959
rect 254667 290931 254701 290959
rect 254729 290931 254763 290959
rect 254791 290931 263577 290959
rect 263605 290931 263639 290959
rect 263667 290931 263701 290959
rect 263729 290931 263763 290959
rect 263791 290931 272577 290959
rect 272605 290931 272639 290959
rect 272667 290931 272701 290959
rect 272729 290931 272763 290959
rect 272791 290931 281577 290959
rect 281605 290931 281639 290959
rect 281667 290931 281701 290959
rect 281729 290931 281763 290959
rect 281791 290931 290577 290959
rect 290605 290931 290639 290959
rect 290667 290931 290701 290959
rect 290729 290931 290763 290959
rect 290791 290931 299256 290959
rect 299284 290931 299318 290959
rect 299346 290931 299380 290959
rect 299408 290931 299442 290959
rect 299470 290931 299998 290959
rect -6 290897 299998 290931
rect -6 290869 522 290897
rect 550 290869 584 290897
rect 612 290869 646 290897
rect 674 290869 708 290897
rect 736 290869 2577 290897
rect 2605 290869 2639 290897
rect 2667 290869 2701 290897
rect 2729 290869 2763 290897
rect 2791 290869 11577 290897
rect 11605 290869 11639 290897
rect 11667 290869 11701 290897
rect 11729 290869 11763 290897
rect 11791 290869 20577 290897
rect 20605 290869 20639 290897
rect 20667 290869 20701 290897
rect 20729 290869 20763 290897
rect 20791 290869 29577 290897
rect 29605 290869 29639 290897
rect 29667 290869 29701 290897
rect 29729 290869 29763 290897
rect 29791 290869 38577 290897
rect 38605 290869 38639 290897
rect 38667 290869 38701 290897
rect 38729 290869 38763 290897
rect 38791 290869 47577 290897
rect 47605 290869 47639 290897
rect 47667 290869 47701 290897
rect 47729 290869 47763 290897
rect 47791 290869 56577 290897
rect 56605 290869 56639 290897
rect 56667 290869 56701 290897
rect 56729 290869 56763 290897
rect 56791 290869 65577 290897
rect 65605 290869 65639 290897
rect 65667 290869 65701 290897
rect 65729 290869 65763 290897
rect 65791 290869 74577 290897
rect 74605 290869 74639 290897
rect 74667 290869 74701 290897
rect 74729 290869 74763 290897
rect 74791 290869 83577 290897
rect 83605 290869 83639 290897
rect 83667 290869 83701 290897
rect 83729 290869 83763 290897
rect 83791 290869 92577 290897
rect 92605 290869 92639 290897
rect 92667 290869 92701 290897
rect 92729 290869 92763 290897
rect 92791 290869 101577 290897
rect 101605 290869 101639 290897
rect 101667 290869 101701 290897
rect 101729 290869 101763 290897
rect 101791 290869 110577 290897
rect 110605 290869 110639 290897
rect 110667 290869 110701 290897
rect 110729 290869 110763 290897
rect 110791 290869 119577 290897
rect 119605 290869 119639 290897
rect 119667 290869 119701 290897
rect 119729 290869 119763 290897
rect 119791 290869 128577 290897
rect 128605 290869 128639 290897
rect 128667 290869 128701 290897
rect 128729 290869 128763 290897
rect 128791 290869 137577 290897
rect 137605 290869 137639 290897
rect 137667 290869 137701 290897
rect 137729 290869 137763 290897
rect 137791 290869 146577 290897
rect 146605 290869 146639 290897
rect 146667 290869 146701 290897
rect 146729 290869 146763 290897
rect 146791 290869 155577 290897
rect 155605 290869 155639 290897
rect 155667 290869 155701 290897
rect 155729 290869 155763 290897
rect 155791 290869 164577 290897
rect 164605 290869 164639 290897
rect 164667 290869 164701 290897
rect 164729 290869 164763 290897
rect 164791 290869 173577 290897
rect 173605 290869 173639 290897
rect 173667 290869 173701 290897
rect 173729 290869 173763 290897
rect 173791 290869 182577 290897
rect 182605 290869 182639 290897
rect 182667 290869 182701 290897
rect 182729 290869 182763 290897
rect 182791 290869 191577 290897
rect 191605 290869 191639 290897
rect 191667 290869 191701 290897
rect 191729 290869 191763 290897
rect 191791 290869 200577 290897
rect 200605 290869 200639 290897
rect 200667 290869 200701 290897
rect 200729 290869 200763 290897
rect 200791 290869 209577 290897
rect 209605 290869 209639 290897
rect 209667 290869 209701 290897
rect 209729 290869 209763 290897
rect 209791 290869 218577 290897
rect 218605 290869 218639 290897
rect 218667 290869 218701 290897
rect 218729 290869 218763 290897
rect 218791 290869 227577 290897
rect 227605 290869 227639 290897
rect 227667 290869 227701 290897
rect 227729 290869 227763 290897
rect 227791 290869 236577 290897
rect 236605 290869 236639 290897
rect 236667 290869 236701 290897
rect 236729 290869 236763 290897
rect 236791 290869 245577 290897
rect 245605 290869 245639 290897
rect 245667 290869 245701 290897
rect 245729 290869 245763 290897
rect 245791 290869 254577 290897
rect 254605 290869 254639 290897
rect 254667 290869 254701 290897
rect 254729 290869 254763 290897
rect 254791 290869 263577 290897
rect 263605 290869 263639 290897
rect 263667 290869 263701 290897
rect 263729 290869 263763 290897
rect 263791 290869 272577 290897
rect 272605 290869 272639 290897
rect 272667 290869 272701 290897
rect 272729 290869 272763 290897
rect 272791 290869 281577 290897
rect 281605 290869 281639 290897
rect 281667 290869 281701 290897
rect 281729 290869 281763 290897
rect 281791 290869 290577 290897
rect 290605 290869 290639 290897
rect 290667 290869 290701 290897
rect 290729 290869 290763 290897
rect 290791 290869 299256 290897
rect 299284 290869 299318 290897
rect 299346 290869 299380 290897
rect 299408 290869 299442 290897
rect 299470 290869 299998 290897
rect -6 290835 299998 290869
rect -6 290807 522 290835
rect 550 290807 584 290835
rect 612 290807 646 290835
rect 674 290807 708 290835
rect 736 290807 2577 290835
rect 2605 290807 2639 290835
rect 2667 290807 2701 290835
rect 2729 290807 2763 290835
rect 2791 290807 11577 290835
rect 11605 290807 11639 290835
rect 11667 290807 11701 290835
rect 11729 290807 11763 290835
rect 11791 290807 20577 290835
rect 20605 290807 20639 290835
rect 20667 290807 20701 290835
rect 20729 290807 20763 290835
rect 20791 290807 29577 290835
rect 29605 290807 29639 290835
rect 29667 290807 29701 290835
rect 29729 290807 29763 290835
rect 29791 290807 38577 290835
rect 38605 290807 38639 290835
rect 38667 290807 38701 290835
rect 38729 290807 38763 290835
rect 38791 290807 47577 290835
rect 47605 290807 47639 290835
rect 47667 290807 47701 290835
rect 47729 290807 47763 290835
rect 47791 290807 56577 290835
rect 56605 290807 56639 290835
rect 56667 290807 56701 290835
rect 56729 290807 56763 290835
rect 56791 290807 65577 290835
rect 65605 290807 65639 290835
rect 65667 290807 65701 290835
rect 65729 290807 65763 290835
rect 65791 290807 74577 290835
rect 74605 290807 74639 290835
rect 74667 290807 74701 290835
rect 74729 290807 74763 290835
rect 74791 290807 83577 290835
rect 83605 290807 83639 290835
rect 83667 290807 83701 290835
rect 83729 290807 83763 290835
rect 83791 290807 92577 290835
rect 92605 290807 92639 290835
rect 92667 290807 92701 290835
rect 92729 290807 92763 290835
rect 92791 290807 101577 290835
rect 101605 290807 101639 290835
rect 101667 290807 101701 290835
rect 101729 290807 101763 290835
rect 101791 290807 110577 290835
rect 110605 290807 110639 290835
rect 110667 290807 110701 290835
rect 110729 290807 110763 290835
rect 110791 290807 119577 290835
rect 119605 290807 119639 290835
rect 119667 290807 119701 290835
rect 119729 290807 119763 290835
rect 119791 290807 128577 290835
rect 128605 290807 128639 290835
rect 128667 290807 128701 290835
rect 128729 290807 128763 290835
rect 128791 290807 137577 290835
rect 137605 290807 137639 290835
rect 137667 290807 137701 290835
rect 137729 290807 137763 290835
rect 137791 290807 146577 290835
rect 146605 290807 146639 290835
rect 146667 290807 146701 290835
rect 146729 290807 146763 290835
rect 146791 290807 155577 290835
rect 155605 290807 155639 290835
rect 155667 290807 155701 290835
rect 155729 290807 155763 290835
rect 155791 290807 164577 290835
rect 164605 290807 164639 290835
rect 164667 290807 164701 290835
rect 164729 290807 164763 290835
rect 164791 290807 173577 290835
rect 173605 290807 173639 290835
rect 173667 290807 173701 290835
rect 173729 290807 173763 290835
rect 173791 290807 182577 290835
rect 182605 290807 182639 290835
rect 182667 290807 182701 290835
rect 182729 290807 182763 290835
rect 182791 290807 191577 290835
rect 191605 290807 191639 290835
rect 191667 290807 191701 290835
rect 191729 290807 191763 290835
rect 191791 290807 200577 290835
rect 200605 290807 200639 290835
rect 200667 290807 200701 290835
rect 200729 290807 200763 290835
rect 200791 290807 209577 290835
rect 209605 290807 209639 290835
rect 209667 290807 209701 290835
rect 209729 290807 209763 290835
rect 209791 290807 218577 290835
rect 218605 290807 218639 290835
rect 218667 290807 218701 290835
rect 218729 290807 218763 290835
rect 218791 290807 227577 290835
rect 227605 290807 227639 290835
rect 227667 290807 227701 290835
rect 227729 290807 227763 290835
rect 227791 290807 236577 290835
rect 236605 290807 236639 290835
rect 236667 290807 236701 290835
rect 236729 290807 236763 290835
rect 236791 290807 245577 290835
rect 245605 290807 245639 290835
rect 245667 290807 245701 290835
rect 245729 290807 245763 290835
rect 245791 290807 254577 290835
rect 254605 290807 254639 290835
rect 254667 290807 254701 290835
rect 254729 290807 254763 290835
rect 254791 290807 263577 290835
rect 263605 290807 263639 290835
rect 263667 290807 263701 290835
rect 263729 290807 263763 290835
rect 263791 290807 272577 290835
rect 272605 290807 272639 290835
rect 272667 290807 272701 290835
rect 272729 290807 272763 290835
rect 272791 290807 281577 290835
rect 281605 290807 281639 290835
rect 281667 290807 281701 290835
rect 281729 290807 281763 290835
rect 281791 290807 290577 290835
rect 290605 290807 290639 290835
rect 290667 290807 290701 290835
rect 290729 290807 290763 290835
rect 290791 290807 299256 290835
rect 299284 290807 299318 290835
rect 299346 290807 299380 290835
rect 299408 290807 299442 290835
rect 299470 290807 299998 290835
rect -6 290773 299998 290807
rect -6 290745 522 290773
rect 550 290745 584 290773
rect 612 290745 646 290773
rect 674 290745 708 290773
rect 736 290745 2577 290773
rect 2605 290745 2639 290773
rect 2667 290745 2701 290773
rect 2729 290745 2763 290773
rect 2791 290745 11577 290773
rect 11605 290745 11639 290773
rect 11667 290745 11701 290773
rect 11729 290745 11763 290773
rect 11791 290745 20577 290773
rect 20605 290745 20639 290773
rect 20667 290745 20701 290773
rect 20729 290745 20763 290773
rect 20791 290745 29577 290773
rect 29605 290745 29639 290773
rect 29667 290745 29701 290773
rect 29729 290745 29763 290773
rect 29791 290745 38577 290773
rect 38605 290745 38639 290773
rect 38667 290745 38701 290773
rect 38729 290745 38763 290773
rect 38791 290745 47577 290773
rect 47605 290745 47639 290773
rect 47667 290745 47701 290773
rect 47729 290745 47763 290773
rect 47791 290745 56577 290773
rect 56605 290745 56639 290773
rect 56667 290745 56701 290773
rect 56729 290745 56763 290773
rect 56791 290745 65577 290773
rect 65605 290745 65639 290773
rect 65667 290745 65701 290773
rect 65729 290745 65763 290773
rect 65791 290745 74577 290773
rect 74605 290745 74639 290773
rect 74667 290745 74701 290773
rect 74729 290745 74763 290773
rect 74791 290745 83577 290773
rect 83605 290745 83639 290773
rect 83667 290745 83701 290773
rect 83729 290745 83763 290773
rect 83791 290745 92577 290773
rect 92605 290745 92639 290773
rect 92667 290745 92701 290773
rect 92729 290745 92763 290773
rect 92791 290745 101577 290773
rect 101605 290745 101639 290773
rect 101667 290745 101701 290773
rect 101729 290745 101763 290773
rect 101791 290745 110577 290773
rect 110605 290745 110639 290773
rect 110667 290745 110701 290773
rect 110729 290745 110763 290773
rect 110791 290745 119577 290773
rect 119605 290745 119639 290773
rect 119667 290745 119701 290773
rect 119729 290745 119763 290773
rect 119791 290745 128577 290773
rect 128605 290745 128639 290773
rect 128667 290745 128701 290773
rect 128729 290745 128763 290773
rect 128791 290745 137577 290773
rect 137605 290745 137639 290773
rect 137667 290745 137701 290773
rect 137729 290745 137763 290773
rect 137791 290745 146577 290773
rect 146605 290745 146639 290773
rect 146667 290745 146701 290773
rect 146729 290745 146763 290773
rect 146791 290745 155577 290773
rect 155605 290745 155639 290773
rect 155667 290745 155701 290773
rect 155729 290745 155763 290773
rect 155791 290745 164577 290773
rect 164605 290745 164639 290773
rect 164667 290745 164701 290773
rect 164729 290745 164763 290773
rect 164791 290745 173577 290773
rect 173605 290745 173639 290773
rect 173667 290745 173701 290773
rect 173729 290745 173763 290773
rect 173791 290745 182577 290773
rect 182605 290745 182639 290773
rect 182667 290745 182701 290773
rect 182729 290745 182763 290773
rect 182791 290745 191577 290773
rect 191605 290745 191639 290773
rect 191667 290745 191701 290773
rect 191729 290745 191763 290773
rect 191791 290745 200577 290773
rect 200605 290745 200639 290773
rect 200667 290745 200701 290773
rect 200729 290745 200763 290773
rect 200791 290745 209577 290773
rect 209605 290745 209639 290773
rect 209667 290745 209701 290773
rect 209729 290745 209763 290773
rect 209791 290745 218577 290773
rect 218605 290745 218639 290773
rect 218667 290745 218701 290773
rect 218729 290745 218763 290773
rect 218791 290745 227577 290773
rect 227605 290745 227639 290773
rect 227667 290745 227701 290773
rect 227729 290745 227763 290773
rect 227791 290745 236577 290773
rect 236605 290745 236639 290773
rect 236667 290745 236701 290773
rect 236729 290745 236763 290773
rect 236791 290745 245577 290773
rect 245605 290745 245639 290773
rect 245667 290745 245701 290773
rect 245729 290745 245763 290773
rect 245791 290745 254577 290773
rect 254605 290745 254639 290773
rect 254667 290745 254701 290773
rect 254729 290745 254763 290773
rect 254791 290745 263577 290773
rect 263605 290745 263639 290773
rect 263667 290745 263701 290773
rect 263729 290745 263763 290773
rect 263791 290745 272577 290773
rect 272605 290745 272639 290773
rect 272667 290745 272701 290773
rect 272729 290745 272763 290773
rect 272791 290745 281577 290773
rect 281605 290745 281639 290773
rect 281667 290745 281701 290773
rect 281729 290745 281763 290773
rect 281791 290745 290577 290773
rect 290605 290745 290639 290773
rect 290667 290745 290701 290773
rect 290729 290745 290763 290773
rect 290791 290745 299256 290773
rect 299284 290745 299318 290773
rect 299346 290745 299380 290773
rect 299408 290745 299442 290773
rect 299470 290745 299998 290773
rect -6 290697 299998 290745
rect -6 284959 299998 285007
rect -6 284931 42 284959
rect 70 284931 104 284959
rect 132 284931 166 284959
rect 194 284931 228 284959
rect 256 284931 4437 284959
rect 4465 284931 4499 284959
rect 4527 284931 4561 284959
rect 4589 284931 4623 284959
rect 4651 284931 13437 284959
rect 13465 284931 13499 284959
rect 13527 284931 13561 284959
rect 13589 284931 13623 284959
rect 13651 284931 22437 284959
rect 22465 284931 22499 284959
rect 22527 284931 22561 284959
rect 22589 284931 22623 284959
rect 22651 284931 31437 284959
rect 31465 284931 31499 284959
rect 31527 284931 31561 284959
rect 31589 284931 31623 284959
rect 31651 284931 40437 284959
rect 40465 284931 40499 284959
rect 40527 284931 40561 284959
rect 40589 284931 40623 284959
rect 40651 284931 49437 284959
rect 49465 284931 49499 284959
rect 49527 284931 49561 284959
rect 49589 284931 49623 284959
rect 49651 284931 58437 284959
rect 58465 284931 58499 284959
rect 58527 284931 58561 284959
rect 58589 284931 58623 284959
rect 58651 284931 67437 284959
rect 67465 284931 67499 284959
rect 67527 284931 67561 284959
rect 67589 284931 67623 284959
rect 67651 284931 76437 284959
rect 76465 284931 76499 284959
rect 76527 284931 76561 284959
rect 76589 284931 76623 284959
rect 76651 284931 85437 284959
rect 85465 284931 85499 284959
rect 85527 284931 85561 284959
rect 85589 284931 85623 284959
rect 85651 284931 94437 284959
rect 94465 284931 94499 284959
rect 94527 284931 94561 284959
rect 94589 284931 94623 284959
rect 94651 284931 103437 284959
rect 103465 284931 103499 284959
rect 103527 284931 103561 284959
rect 103589 284931 103623 284959
rect 103651 284931 112437 284959
rect 112465 284931 112499 284959
rect 112527 284931 112561 284959
rect 112589 284931 112623 284959
rect 112651 284931 121437 284959
rect 121465 284931 121499 284959
rect 121527 284931 121561 284959
rect 121589 284931 121623 284959
rect 121651 284931 130437 284959
rect 130465 284931 130499 284959
rect 130527 284931 130561 284959
rect 130589 284931 130623 284959
rect 130651 284931 139437 284959
rect 139465 284931 139499 284959
rect 139527 284931 139561 284959
rect 139589 284931 139623 284959
rect 139651 284931 148437 284959
rect 148465 284931 148499 284959
rect 148527 284931 148561 284959
rect 148589 284931 148623 284959
rect 148651 284931 157437 284959
rect 157465 284931 157499 284959
rect 157527 284931 157561 284959
rect 157589 284931 157623 284959
rect 157651 284931 166437 284959
rect 166465 284931 166499 284959
rect 166527 284931 166561 284959
rect 166589 284931 166623 284959
rect 166651 284931 175437 284959
rect 175465 284931 175499 284959
rect 175527 284931 175561 284959
rect 175589 284931 175623 284959
rect 175651 284931 184437 284959
rect 184465 284931 184499 284959
rect 184527 284931 184561 284959
rect 184589 284931 184623 284959
rect 184651 284931 193437 284959
rect 193465 284931 193499 284959
rect 193527 284931 193561 284959
rect 193589 284931 193623 284959
rect 193651 284931 202437 284959
rect 202465 284931 202499 284959
rect 202527 284931 202561 284959
rect 202589 284931 202623 284959
rect 202651 284931 211437 284959
rect 211465 284931 211499 284959
rect 211527 284931 211561 284959
rect 211589 284931 211623 284959
rect 211651 284931 220437 284959
rect 220465 284931 220499 284959
rect 220527 284931 220561 284959
rect 220589 284931 220623 284959
rect 220651 284931 229437 284959
rect 229465 284931 229499 284959
rect 229527 284931 229561 284959
rect 229589 284931 229623 284959
rect 229651 284931 238437 284959
rect 238465 284931 238499 284959
rect 238527 284931 238561 284959
rect 238589 284931 238623 284959
rect 238651 284931 247437 284959
rect 247465 284931 247499 284959
rect 247527 284931 247561 284959
rect 247589 284931 247623 284959
rect 247651 284931 256437 284959
rect 256465 284931 256499 284959
rect 256527 284931 256561 284959
rect 256589 284931 256623 284959
rect 256651 284931 265437 284959
rect 265465 284931 265499 284959
rect 265527 284931 265561 284959
rect 265589 284931 265623 284959
rect 265651 284931 274437 284959
rect 274465 284931 274499 284959
rect 274527 284931 274561 284959
rect 274589 284931 274623 284959
rect 274651 284931 283437 284959
rect 283465 284931 283499 284959
rect 283527 284931 283561 284959
rect 283589 284931 283623 284959
rect 283651 284931 292437 284959
rect 292465 284931 292499 284959
rect 292527 284931 292561 284959
rect 292589 284931 292623 284959
rect 292651 284931 299736 284959
rect 299764 284931 299798 284959
rect 299826 284931 299860 284959
rect 299888 284931 299922 284959
rect 299950 284931 299998 284959
rect -6 284897 299998 284931
rect -6 284869 42 284897
rect 70 284869 104 284897
rect 132 284869 166 284897
rect 194 284869 228 284897
rect 256 284869 4437 284897
rect 4465 284869 4499 284897
rect 4527 284869 4561 284897
rect 4589 284869 4623 284897
rect 4651 284869 13437 284897
rect 13465 284869 13499 284897
rect 13527 284869 13561 284897
rect 13589 284869 13623 284897
rect 13651 284869 22437 284897
rect 22465 284869 22499 284897
rect 22527 284869 22561 284897
rect 22589 284869 22623 284897
rect 22651 284869 31437 284897
rect 31465 284869 31499 284897
rect 31527 284869 31561 284897
rect 31589 284869 31623 284897
rect 31651 284869 40437 284897
rect 40465 284869 40499 284897
rect 40527 284869 40561 284897
rect 40589 284869 40623 284897
rect 40651 284869 49437 284897
rect 49465 284869 49499 284897
rect 49527 284869 49561 284897
rect 49589 284869 49623 284897
rect 49651 284869 58437 284897
rect 58465 284869 58499 284897
rect 58527 284869 58561 284897
rect 58589 284869 58623 284897
rect 58651 284869 67437 284897
rect 67465 284869 67499 284897
rect 67527 284869 67561 284897
rect 67589 284869 67623 284897
rect 67651 284869 76437 284897
rect 76465 284869 76499 284897
rect 76527 284869 76561 284897
rect 76589 284869 76623 284897
rect 76651 284869 85437 284897
rect 85465 284869 85499 284897
rect 85527 284869 85561 284897
rect 85589 284869 85623 284897
rect 85651 284869 94437 284897
rect 94465 284869 94499 284897
rect 94527 284869 94561 284897
rect 94589 284869 94623 284897
rect 94651 284869 103437 284897
rect 103465 284869 103499 284897
rect 103527 284869 103561 284897
rect 103589 284869 103623 284897
rect 103651 284869 112437 284897
rect 112465 284869 112499 284897
rect 112527 284869 112561 284897
rect 112589 284869 112623 284897
rect 112651 284869 121437 284897
rect 121465 284869 121499 284897
rect 121527 284869 121561 284897
rect 121589 284869 121623 284897
rect 121651 284869 130437 284897
rect 130465 284869 130499 284897
rect 130527 284869 130561 284897
rect 130589 284869 130623 284897
rect 130651 284869 139437 284897
rect 139465 284869 139499 284897
rect 139527 284869 139561 284897
rect 139589 284869 139623 284897
rect 139651 284869 148437 284897
rect 148465 284869 148499 284897
rect 148527 284869 148561 284897
rect 148589 284869 148623 284897
rect 148651 284869 157437 284897
rect 157465 284869 157499 284897
rect 157527 284869 157561 284897
rect 157589 284869 157623 284897
rect 157651 284869 166437 284897
rect 166465 284869 166499 284897
rect 166527 284869 166561 284897
rect 166589 284869 166623 284897
rect 166651 284869 175437 284897
rect 175465 284869 175499 284897
rect 175527 284869 175561 284897
rect 175589 284869 175623 284897
rect 175651 284869 184437 284897
rect 184465 284869 184499 284897
rect 184527 284869 184561 284897
rect 184589 284869 184623 284897
rect 184651 284869 193437 284897
rect 193465 284869 193499 284897
rect 193527 284869 193561 284897
rect 193589 284869 193623 284897
rect 193651 284869 202437 284897
rect 202465 284869 202499 284897
rect 202527 284869 202561 284897
rect 202589 284869 202623 284897
rect 202651 284869 211437 284897
rect 211465 284869 211499 284897
rect 211527 284869 211561 284897
rect 211589 284869 211623 284897
rect 211651 284869 220437 284897
rect 220465 284869 220499 284897
rect 220527 284869 220561 284897
rect 220589 284869 220623 284897
rect 220651 284869 229437 284897
rect 229465 284869 229499 284897
rect 229527 284869 229561 284897
rect 229589 284869 229623 284897
rect 229651 284869 238437 284897
rect 238465 284869 238499 284897
rect 238527 284869 238561 284897
rect 238589 284869 238623 284897
rect 238651 284869 247437 284897
rect 247465 284869 247499 284897
rect 247527 284869 247561 284897
rect 247589 284869 247623 284897
rect 247651 284869 256437 284897
rect 256465 284869 256499 284897
rect 256527 284869 256561 284897
rect 256589 284869 256623 284897
rect 256651 284869 265437 284897
rect 265465 284869 265499 284897
rect 265527 284869 265561 284897
rect 265589 284869 265623 284897
rect 265651 284869 274437 284897
rect 274465 284869 274499 284897
rect 274527 284869 274561 284897
rect 274589 284869 274623 284897
rect 274651 284869 283437 284897
rect 283465 284869 283499 284897
rect 283527 284869 283561 284897
rect 283589 284869 283623 284897
rect 283651 284869 292437 284897
rect 292465 284869 292499 284897
rect 292527 284869 292561 284897
rect 292589 284869 292623 284897
rect 292651 284869 299736 284897
rect 299764 284869 299798 284897
rect 299826 284869 299860 284897
rect 299888 284869 299922 284897
rect 299950 284869 299998 284897
rect -6 284835 299998 284869
rect -6 284807 42 284835
rect 70 284807 104 284835
rect 132 284807 166 284835
rect 194 284807 228 284835
rect 256 284807 4437 284835
rect 4465 284807 4499 284835
rect 4527 284807 4561 284835
rect 4589 284807 4623 284835
rect 4651 284807 13437 284835
rect 13465 284807 13499 284835
rect 13527 284807 13561 284835
rect 13589 284807 13623 284835
rect 13651 284807 22437 284835
rect 22465 284807 22499 284835
rect 22527 284807 22561 284835
rect 22589 284807 22623 284835
rect 22651 284807 31437 284835
rect 31465 284807 31499 284835
rect 31527 284807 31561 284835
rect 31589 284807 31623 284835
rect 31651 284807 40437 284835
rect 40465 284807 40499 284835
rect 40527 284807 40561 284835
rect 40589 284807 40623 284835
rect 40651 284807 49437 284835
rect 49465 284807 49499 284835
rect 49527 284807 49561 284835
rect 49589 284807 49623 284835
rect 49651 284807 58437 284835
rect 58465 284807 58499 284835
rect 58527 284807 58561 284835
rect 58589 284807 58623 284835
rect 58651 284807 67437 284835
rect 67465 284807 67499 284835
rect 67527 284807 67561 284835
rect 67589 284807 67623 284835
rect 67651 284807 76437 284835
rect 76465 284807 76499 284835
rect 76527 284807 76561 284835
rect 76589 284807 76623 284835
rect 76651 284807 85437 284835
rect 85465 284807 85499 284835
rect 85527 284807 85561 284835
rect 85589 284807 85623 284835
rect 85651 284807 94437 284835
rect 94465 284807 94499 284835
rect 94527 284807 94561 284835
rect 94589 284807 94623 284835
rect 94651 284807 103437 284835
rect 103465 284807 103499 284835
rect 103527 284807 103561 284835
rect 103589 284807 103623 284835
rect 103651 284807 112437 284835
rect 112465 284807 112499 284835
rect 112527 284807 112561 284835
rect 112589 284807 112623 284835
rect 112651 284807 121437 284835
rect 121465 284807 121499 284835
rect 121527 284807 121561 284835
rect 121589 284807 121623 284835
rect 121651 284807 130437 284835
rect 130465 284807 130499 284835
rect 130527 284807 130561 284835
rect 130589 284807 130623 284835
rect 130651 284807 139437 284835
rect 139465 284807 139499 284835
rect 139527 284807 139561 284835
rect 139589 284807 139623 284835
rect 139651 284807 148437 284835
rect 148465 284807 148499 284835
rect 148527 284807 148561 284835
rect 148589 284807 148623 284835
rect 148651 284807 157437 284835
rect 157465 284807 157499 284835
rect 157527 284807 157561 284835
rect 157589 284807 157623 284835
rect 157651 284807 166437 284835
rect 166465 284807 166499 284835
rect 166527 284807 166561 284835
rect 166589 284807 166623 284835
rect 166651 284807 175437 284835
rect 175465 284807 175499 284835
rect 175527 284807 175561 284835
rect 175589 284807 175623 284835
rect 175651 284807 184437 284835
rect 184465 284807 184499 284835
rect 184527 284807 184561 284835
rect 184589 284807 184623 284835
rect 184651 284807 193437 284835
rect 193465 284807 193499 284835
rect 193527 284807 193561 284835
rect 193589 284807 193623 284835
rect 193651 284807 202437 284835
rect 202465 284807 202499 284835
rect 202527 284807 202561 284835
rect 202589 284807 202623 284835
rect 202651 284807 211437 284835
rect 211465 284807 211499 284835
rect 211527 284807 211561 284835
rect 211589 284807 211623 284835
rect 211651 284807 220437 284835
rect 220465 284807 220499 284835
rect 220527 284807 220561 284835
rect 220589 284807 220623 284835
rect 220651 284807 229437 284835
rect 229465 284807 229499 284835
rect 229527 284807 229561 284835
rect 229589 284807 229623 284835
rect 229651 284807 238437 284835
rect 238465 284807 238499 284835
rect 238527 284807 238561 284835
rect 238589 284807 238623 284835
rect 238651 284807 247437 284835
rect 247465 284807 247499 284835
rect 247527 284807 247561 284835
rect 247589 284807 247623 284835
rect 247651 284807 256437 284835
rect 256465 284807 256499 284835
rect 256527 284807 256561 284835
rect 256589 284807 256623 284835
rect 256651 284807 265437 284835
rect 265465 284807 265499 284835
rect 265527 284807 265561 284835
rect 265589 284807 265623 284835
rect 265651 284807 274437 284835
rect 274465 284807 274499 284835
rect 274527 284807 274561 284835
rect 274589 284807 274623 284835
rect 274651 284807 283437 284835
rect 283465 284807 283499 284835
rect 283527 284807 283561 284835
rect 283589 284807 283623 284835
rect 283651 284807 292437 284835
rect 292465 284807 292499 284835
rect 292527 284807 292561 284835
rect 292589 284807 292623 284835
rect 292651 284807 299736 284835
rect 299764 284807 299798 284835
rect 299826 284807 299860 284835
rect 299888 284807 299922 284835
rect 299950 284807 299998 284835
rect -6 284773 299998 284807
rect -6 284745 42 284773
rect 70 284745 104 284773
rect 132 284745 166 284773
rect 194 284745 228 284773
rect 256 284745 4437 284773
rect 4465 284745 4499 284773
rect 4527 284745 4561 284773
rect 4589 284745 4623 284773
rect 4651 284745 13437 284773
rect 13465 284745 13499 284773
rect 13527 284745 13561 284773
rect 13589 284745 13623 284773
rect 13651 284745 22437 284773
rect 22465 284745 22499 284773
rect 22527 284745 22561 284773
rect 22589 284745 22623 284773
rect 22651 284745 31437 284773
rect 31465 284745 31499 284773
rect 31527 284745 31561 284773
rect 31589 284745 31623 284773
rect 31651 284745 40437 284773
rect 40465 284745 40499 284773
rect 40527 284745 40561 284773
rect 40589 284745 40623 284773
rect 40651 284745 49437 284773
rect 49465 284745 49499 284773
rect 49527 284745 49561 284773
rect 49589 284745 49623 284773
rect 49651 284745 58437 284773
rect 58465 284745 58499 284773
rect 58527 284745 58561 284773
rect 58589 284745 58623 284773
rect 58651 284745 67437 284773
rect 67465 284745 67499 284773
rect 67527 284745 67561 284773
rect 67589 284745 67623 284773
rect 67651 284745 76437 284773
rect 76465 284745 76499 284773
rect 76527 284745 76561 284773
rect 76589 284745 76623 284773
rect 76651 284745 85437 284773
rect 85465 284745 85499 284773
rect 85527 284745 85561 284773
rect 85589 284745 85623 284773
rect 85651 284745 94437 284773
rect 94465 284745 94499 284773
rect 94527 284745 94561 284773
rect 94589 284745 94623 284773
rect 94651 284745 103437 284773
rect 103465 284745 103499 284773
rect 103527 284745 103561 284773
rect 103589 284745 103623 284773
rect 103651 284745 112437 284773
rect 112465 284745 112499 284773
rect 112527 284745 112561 284773
rect 112589 284745 112623 284773
rect 112651 284745 121437 284773
rect 121465 284745 121499 284773
rect 121527 284745 121561 284773
rect 121589 284745 121623 284773
rect 121651 284745 130437 284773
rect 130465 284745 130499 284773
rect 130527 284745 130561 284773
rect 130589 284745 130623 284773
rect 130651 284745 139437 284773
rect 139465 284745 139499 284773
rect 139527 284745 139561 284773
rect 139589 284745 139623 284773
rect 139651 284745 148437 284773
rect 148465 284745 148499 284773
rect 148527 284745 148561 284773
rect 148589 284745 148623 284773
rect 148651 284745 157437 284773
rect 157465 284745 157499 284773
rect 157527 284745 157561 284773
rect 157589 284745 157623 284773
rect 157651 284745 166437 284773
rect 166465 284745 166499 284773
rect 166527 284745 166561 284773
rect 166589 284745 166623 284773
rect 166651 284745 175437 284773
rect 175465 284745 175499 284773
rect 175527 284745 175561 284773
rect 175589 284745 175623 284773
rect 175651 284745 184437 284773
rect 184465 284745 184499 284773
rect 184527 284745 184561 284773
rect 184589 284745 184623 284773
rect 184651 284745 193437 284773
rect 193465 284745 193499 284773
rect 193527 284745 193561 284773
rect 193589 284745 193623 284773
rect 193651 284745 202437 284773
rect 202465 284745 202499 284773
rect 202527 284745 202561 284773
rect 202589 284745 202623 284773
rect 202651 284745 211437 284773
rect 211465 284745 211499 284773
rect 211527 284745 211561 284773
rect 211589 284745 211623 284773
rect 211651 284745 220437 284773
rect 220465 284745 220499 284773
rect 220527 284745 220561 284773
rect 220589 284745 220623 284773
rect 220651 284745 229437 284773
rect 229465 284745 229499 284773
rect 229527 284745 229561 284773
rect 229589 284745 229623 284773
rect 229651 284745 238437 284773
rect 238465 284745 238499 284773
rect 238527 284745 238561 284773
rect 238589 284745 238623 284773
rect 238651 284745 247437 284773
rect 247465 284745 247499 284773
rect 247527 284745 247561 284773
rect 247589 284745 247623 284773
rect 247651 284745 256437 284773
rect 256465 284745 256499 284773
rect 256527 284745 256561 284773
rect 256589 284745 256623 284773
rect 256651 284745 265437 284773
rect 265465 284745 265499 284773
rect 265527 284745 265561 284773
rect 265589 284745 265623 284773
rect 265651 284745 274437 284773
rect 274465 284745 274499 284773
rect 274527 284745 274561 284773
rect 274589 284745 274623 284773
rect 274651 284745 283437 284773
rect 283465 284745 283499 284773
rect 283527 284745 283561 284773
rect 283589 284745 283623 284773
rect 283651 284745 292437 284773
rect 292465 284745 292499 284773
rect 292527 284745 292561 284773
rect 292589 284745 292623 284773
rect 292651 284745 299736 284773
rect 299764 284745 299798 284773
rect 299826 284745 299860 284773
rect 299888 284745 299922 284773
rect 299950 284745 299998 284773
rect -6 284697 299998 284745
rect -6 281959 299998 282007
rect -6 281931 522 281959
rect 550 281931 584 281959
rect 612 281931 646 281959
rect 674 281931 708 281959
rect 736 281931 2577 281959
rect 2605 281931 2639 281959
rect 2667 281931 2701 281959
rect 2729 281931 2763 281959
rect 2791 281931 11577 281959
rect 11605 281931 11639 281959
rect 11667 281931 11701 281959
rect 11729 281931 11763 281959
rect 11791 281931 20577 281959
rect 20605 281931 20639 281959
rect 20667 281931 20701 281959
rect 20729 281931 20763 281959
rect 20791 281931 29577 281959
rect 29605 281931 29639 281959
rect 29667 281931 29701 281959
rect 29729 281931 29763 281959
rect 29791 281931 38577 281959
rect 38605 281931 38639 281959
rect 38667 281931 38701 281959
rect 38729 281931 38763 281959
rect 38791 281931 47577 281959
rect 47605 281931 47639 281959
rect 47667 281931 47701 281959
rect 47729 281931 47763 281959
rect 47791 281931 56577 281959
rect 56605 281931 56639 281959
rect 56667 281931 56701 281959
rect 56729 281931 56763 281959
rect 56791 281931 65577 281959
rect 65605 281931 65639 281959
rect 65667 281931 65701 281959
rect 65729 281931 65763 281959
rect 65791 281931 74577 281959
rect 74605 281931 74639 281959
rect 74667 281931 74701 281959
rect 74729 281931 74763 281959
rect 74791 281931 83577 281959
rect 83605 281931 83639 281959
rect 83667 281931 83701 281959
rect 83729 281931 83763 281959
rect 83791 281931 92577 281959
rect 92605 281931 92639 281959
rect 92667 281931 92701 281959
rect 92729 281931 92763 281959
rect 92791 281931 101577 281959
rect 101605 281931 101639 281959
rect 101667 281931 101701 281959
rect 101729 281931 101763 281959
rect 101791 281931 110577 281959
rect 110605 281931 110639 281959
rect 110667 281931 110701 281959
rect 110729 281931 110763 281959
rect 110791 281931 119577 281959
rect 119605 281931 119639 281959
rect 119667 281931 119701 281959
rect 119729 281931 119763 281959
rect 119791 281931 128577 281959
rect 128605 281931 128639 281959
rect 128667 281931 128701 281959
rect 128729 281931 128763 281959
rect 128791 281931 137577 281959
rect 137605 281931 137639 281959
rect 137667 281931 137701 281959
rect 137729 281931 137763 281959
rect 137791 281931 146577 281959
rect 146605 281931 146639 281959
rect 146667 281931 146701 281959
rect 146729 281931 146763 281959
rect 146791 281931 155577 281959
rect 155605 281931 155639 281959
rect 155667 281931 155701 281959
rect 155729 281931 155763 281959
rect 155791 281931 164577 281959
rect 164605 281931 164639 281959
rect 164667 281931 164701 281959
rect 164729 281931 164763 281959
rect 164791 281931 173577 281959
rect 173605 281931 173639 281959
rect 173667 281931 173701 281959
rect 173729 281931 173763 281959
rect 173791 281931 182577 281959
rect 182605 281931 182639 281959
rect 182667 281931 182701 281959
rect 182729 281931 182763 281959
rect 182791 281931 191577 281959
rect 191605 281931 191639 281959
rect 191667 281931 191701 281959
rect 191729 281931 191763 281959
rect 191791 281931 200577 281959
rect 200605 281931 200639 281959
rect 200667 281931 200701 281959
rect 200729 281931 200763 281959
rect 200791 281931 209577 281959
rect 209605 281931 209639 281959
rect 209667 281931 209701 281959
rect 209729 281931 209763 281959
rect 209791 281931 218577 281959
rect 218605 281931 218639 281959
rect 218667 281931 218701 281959
rect 218729 281931 218763 281959
rect 218791 281931 227577 281959
rect 227605 281931 227639 281959
rect 227667 281931 227701 281959
rect 227729 281931 227763 281959
rect 227791 281931 236577 281959
rect 236605 281931 236639 281959
rect 236667 281931 236701 281959
rect 236729 281931 236763 281959
rect 236791 281931 245577 281959
rect 245605 281931 245639 281959
rect 245667 281931 245701 281959
rect 245729 281931 245763 281959
rect 245791 281931 254577 281959
rect 254605 281931 254639 281959
rect 254667 281931 254701 281959
rect 254729 281931 254763 281959
rect 254791 281931 263577 281959
rect 263605 281931 263639 281959
rect 263667 281931 263701 281959
rect 263729 281931 263763 281959
rect 263791 281931 272577 281959
rect 272605 281931 272639 281959
rect 272667 281931 272701 281959
rect 272729 281931 272763 281959
rect 272791 281931 281577 281959
rect 281605 281931 281639 281959
rect 281667 281931 281701 281959
rect 281729 281931 281763 281959
rect 281791 281931 290577 281959
rect 290605 281931 290639 281959
rect 290667 281931 290701 281959
rect 290729 281931 290763 281959
rect 290791 281931 299256 281959
rect 299284 281931 299318 281959
rect 299346 281931 299380 281959
rect 299408 281931 299442 281959
rect 299470 281931 299998 281959
rect -6 281897 299998 281931
rect -6 281869 522 281897
rect 550 281869 584 281897
rect 612 281869 646 281897
rect 674 281869 708 281897
rect 736 281869 2577 281897
rect 2605 281869 2639 281897
rect 2667 281869 2701 281897
rect 2729 281869 2763 281897
rect 2791 281869 11577 281897
rect 11605 281869 11639 281897
rect 11667 281869 11701 281897
rect 11729 281869 11763 281897
rect 11791 281869 20577 281897
rect 20605 281869 20639 281897
rect 20667 281869 20701 281897
rect 20729 281869 20763 281897
rect 20791 281869 29577 281897
rect 29605 281869 29639 281897
rect 29667 281869 29701 281897
rect 29729 281869 29763 281897
rect 29791 281869 38577 281897
rect 38605 281869 38639 281897
rect 38667 281869 38701 281897
rect 38729 281869 38763 281897
rect 38791 281869 47577 281897
rect 47605 281869 47639 281897
rect 47667 281869 47701 281897
rect 47729 281869 47763 281897
rect 47791 281869 56577 281897
rect 56605 281869 56639 281897
rect 56667 281869 56701 281897
rect 56729 281869 56763 281897
rect 56791 281869 65577 281897
rect 65605 281869 65639 281897
rect 65667 281869 65701 281897
rect 65729 281869 65763 281897
rect 65791 281869 74577 281897
rect 74605 281869 74639 281897
rect 74667 281869 74701 281897
rect 74729 281869 74763 281897
rect 74791 281869 83577 281897
rect 83605 281869 83639 281897
rect 83667 281869 83701 281897
rect 83729 281869 83763 281897
rect 83791 281869 92577 281897
rect 92605 281869 92639 281897
rect 92667 281869 92701 281897
rect 92729 281869 92763 281897
rect 92791 281869 101577 281897
rect 101605 281869 101639 281897
rect 101667 281869 101701 281897
rect 101729 281869 101763 281897
rect 101791 281869 110577 281897
rect 110605 281869 110639 281897
rect 110667 281869 110701 281897
rect 110729 281869 110763 281897
rect 110791 281869 119577 281897
rect 119605 281869 119639 281897
rect 119667 281869 119701 281897
rect 119729 281869 119763 281897
rect 119791 281869 128577 281897
rect 128605 281869 128639 281897
rect 128667 281869 128701 281897
rect 128729 281869 128763 281897
rect 128791 281869 137577 281897
rect 137605 281869 137639 281897
rect 137667 281869 137701 281897
rect 137729 281869 137763 281897
rect 137791 281869 146577 281897
rect 146605 281869 146639 281897
rect 146667 281869 146701 281897
rect 146729 281869 146763 281897
rect 146791 281869 155577 281897
rect 155605 281869 155639 281897
rect 155667 281869 155701 281897
rect 155729 281869 155763 281897
rect 155791 281869 164577 281897
rect 164605 281869 164639 281897
rect 164667 281869 164701 281897
rect 164729 281869 164763 281897
rect 164791 281869 173577 281897
rect 173605 281869 173639 281897
rect 173667 281869 173701 281897
rect 173729 281869 173763 281897
rect 173791 281869 182577 281897
rect 182605 281869 182639 281897
rect 182667 281869 182701 281897
rect 182729 281869 182763 281897
rect 182791 281869 191577 281897
rect 191605 281869 191639 281897
rect 191667 281869 191701 281897
rect 191729 281869 191763 281897
rect 191791 281869 200577 281897
rect 200605 281869 200639 281897
rect 200667 281869 200701 281897
rect 200729 281869 200763 281897
rect 200791 281869 209577 281897
rect 209605 281869 209639 281897
rect 209667 281869 209701 281897
rect 209729 281869 209763 281897
rect 209791 281869 218577 281897
rect 218605 281869 218639 281897
rect 218667 281869 218701 281897
rect 218729 281869 218763 281897
rect 218791 281869 227577 281897
rect 227605 281869 227639 281897
rect 227667 281869 227701 281897
rect 227729 281869 227763 281897
rect 227791 281869 236577 281897
rect 236605 281869 236639 281897
rect 236667 281869 236701 281897
rect 236729 281869 236763 281897
rect 236791 281869 245577 281897
rect 245605 281869 245639 281897
rect 245667 281869 245701 281897
rect 245729 281869 245763 281897
rect 245791 281869 254577 281897
rect 254605 281869 254639 281897
rect 254667 281869 254701 281897
rect 254729 281869 254763 281897
rect 254791 281869 263577 281897
rect 263605 281869 263639 281897
rect 263667 281869 263701 281897
rect 263729 281869 263763 281897
rect 263791 281869 272577 281897
rect 272605 281869 272639 281897
rect 272667 281869 272701 281897
rect 272729 281869 272763 281897
rect 272791 281869 281577 281897
rect 281605 281869 281639 281897
rect 281667 281869 281701 281897
rect 281729 281869 281763 281897
rect 281791 281869 290577 281897
rect 290605 281869 290639 281897
rect 290667 281869 290701 281897
rect 290729 281869 290763 281897
rect 290791 281869 299256 281897
rect 299284 281869 299318 281897
rect 299346 281869 299380 281897
rect 299408 281869 299442 281897
rect 299470 281869 299998 281897
rect -6 281835 299998 281869
rect -6 281807 522 281835
rect 550 281807 584 281835
rect 612 281807 646 281835
rect 674 281807 708 281835
rect 736 281807 2577 281835
rect 2605 281807 2639 281835
rect 2667 281807 2701 281835
rect 2729 281807 2763 281835
rect 2791 281807 11577 281835
rect 11605 281807 11639 281835
rect 11667 281807 11701 281835
rect 11729 281807 11763 281835
rect 11791 281807 20577 281835
rect 20605 281807 20639 281835
rect 20667 281807 20701 281835
rect 20729 281807 20763 281835
rect 20791 281807 29577 281835
rect 29605 281807 29639 281835
rect 29667 281807 29701 281835
rect 29729 281807 29763 281835
rect 29791 281807 38577 281835
rect 38605 281807 38639 281835
rect 38667 281807 38701 281835
rect 38729 281807 38763 281835
rect 38791 281807 47577 281835
rect 47605 281807 47639 281835
rect 47667 281807 47701 281835
rect 47729 281807 47763 281835
rect 47791 281807 56577 281835
rect 56605 281807 56639 281835
rect 56667 281807 56701 281835
rect 56729 281807 56763 281835
rect 56791 281807 65577 281835
rect 65605 281807 65639 281835
rect 65667 281807 65701 281835
rect 65729 281807 65763 281835
rect 65791 281807 74577 281835
rect 74605 281807 74639 281835
rect 74667 281807 74701 281835
rect 74729 281807 74763 281835
rect 74791 281807 83577 281835
rect 83605 281807 83639 281835
rect 83667 281807 83701 281835
rect 83729 281807 83763 281835
rect 83791 281807 92577 281835
rect 92605 281807 92639 281835
rect 92667 281807 92701 281835
rect 92729 281807 92763 281835
rect 92791 281807 101577 281835
rect 101605 281807 101639 281835
rect 101667 281807 101701 281835
rect 101729 281807 101763 281835
rect 101791 281807 110577 281835
rect 110605 281807 110639 281835
rect 110667 281807 110701 281835
rect 110729 281807 110763 281835
rect 110791 281807 119577 281835
rect 119605 281807 119639 281835
rect 119667 281807 119701 281835
rect 119729 281807 119763 281835
rect 119791 281807 128577 281835
rect 128605 281807 128639 281835
rect 128667 281807 128701 281835
rect 128729 281807 128763 281835
rect 128791 281807 137577 281835
rect 137605 281807 137639 281835
rect 137667 281807 137701 281835
rect 137729 281807 137763 281835
rect 137791 281807 146577 281835
rect 146605 281807 146639 281835
rect 146667 281807 146701 281835
rect 146729 281807 146763 281835
rect 146791 281807 155577 281835
rect 155605 281807 155639 281835
rect 155667 281807 155701 281835
rect 155729 281807 155763 281835
rect 155791 281807 164577 281835
rect 164605 281807 164639 281835
rect 164667 281807 164701 281835
rect 164729 281807 164763 281835
rect 164791 281807 173577 281835
rect 173605 281807 173639 281835
rect 173667 281807 173701 281835
rect 173729 281807 173763 281835
rect 173791 281807 182577 281835
rect 182605 281807 182639 281835
rect 182667 281807 182701 281835
rect 182729 281807 182763 281835
rect 182791 281807 191577 281835
rect 191605 281807 191639 281835
rect 191667 281807 191701 281835
rect 191729 281807 191763 281835
rect 191791 281807 200577 281835
rect 200605 281807 200639 281835
rect 200667 281807 200701 281835
rect 200729 281807 200763 281835
rect 200791 281807 209577 281835
rect 209605 281807 209639 281835
rect 209667 281807 209701 281835
rect 209729 281807 209763 281835
rect 209791 281807 218577 281835
rect 218605 281807 218639 281835
rect 218667 281807 218701 281835
rect 218729 281807 218763 281835
rect 218791 281807 227577 281835
rect 227605 281807 227639 281835
rect 227667 281807 227701 281835
rect 227729 281807 227763 281835
rect 227791 281807 236577 281835
rect 236605 281807 236639 281835
rect 236667 281807 236701 281835
rect 236729 281807 236763 281835
rect 236791 281807 245577 281835
rect 245605 281807 245639 281835
rect 245667 281807 245701 281835
rect 245729 281807 245763 281835
rect 245791 281807 254577 281835
rect 254605 281807 254639 281835
rect 254667 281807 254701 281835
rect 254729 281807 254763 281835
rect 254791 281807 263577 281835
rect 263605 281807 263639 281835
rect 263667 281807 263701 281835
rect 263729 281807 263763 281835
rect 263791 281807 272577 281835
rect 272605 281807 272639 281835
rect 272667 281807 272701 281835
rect 272729 281807 272763 281835
rect 272791 281807 281577 281835
rect 281605 281807 281639 281835
rect 281667 281807 281701 281835
rect 281729 281807 281763 281835
rect 281791 281807 290577 281835
rect 290605 281807 290639 281835
rect 290667 281807 290701 281835
rect 290729 281807 290763 281835
rect 290791 281807 299256 281835
rect 299284 281807 299318 281835
rect 299346 281807 299380 281835
rect 299408 281807 299442 281835
rect 299470 281807 299998 281835
rect -6 281773 299998 281807
rect -6 281745 522 281773
rect 550 281745 584 281773
rect 612 281745 646 281773
rect 674 281745 708 281773
rect 736 281745 2577 281773
rect 2605 281745 2639 281773
rect 2667 281745 2701 281773
rect 2729 281745 2763 281773
rect 2791 281745 11577 281773
rect 11605 281745 11639 281773
rect 11667 281745 11701 281773
rect 11729 281745 11763 281773
rect 11791 281745 20577 281773
rect 20605 281745 20639 281773
rect 20667 281745 20701 281773
rect 20729 281745 20763 281773
rect 20791 281745 29577 281773
rect 29605 281745 29639 281773
rect 29667 281745 29701 281773
rect 29729 281745 29763 281773
rect 29791 281745 38577 281773
rect 38605 281745 38639 281773
rect 38667 281745 38701 281773
rect 38729 281745 38763 281773
rect 38791 281745 47577 281773
rect 47605 281745 47639 281773
rect 47667 281745 47701 281773
rect 47729 281745 47763 281773
rect 47791 281745 56577 281773
rect 56605 281745 56639 281773
rect 56667 281745 56701 281773
rect 56729 281745 56763 281773
rect 56791 281745 65577 281773
rect 65605 281745 65639 281773
rect 65667 281745 65701 281773
rect 65729 281745 65763 281773
rect 65791 281745 74577 281773
rect 74605 281745 74639 281773
rect 74667 281745 74701 281773
rect 74729 281745 74763 281773
rect 74791 281745 83577 281773
rect 83605 281745 83639 281773
rect 83667 281745 83701 281773
rect 83729 281745 83763 281773
rect 83791 281745 92577 281773
rect 92605 281745 92639 281773
rect 92667 281745 92701 281773
rect 92729 281745 92763 281773
rect 92791 281745 101577 281773
rect 101605 281745 101639 281773
rect 101667 281745 101701 281773
rect 101729 281745 101763 281773
rect 101791 281745 110577 281773
rect 110605 281745 110639 281773
rect 110667 281745 110701 281773
rect 110729 281745 110763 281773
rect 110791 281745 119577 281773
rect 119605 281745 119639 281773
rect 119667 281745 119701 281773
rect 119729 281745 119763 281773
rect 119791 281745 128577 281773
rect 128605 281745 128639 281773
rect 128667 281745 128701 281773
rect 128729 281745 128763 281773
rect 128791 281745 137577 281773
rect 137605 281745 137639 281773
rect 137667 281745 137701 281773
rect 137729 281745 137763 281773
rect 137791 281745 146577 281773
rect 146605 281745 146639 281773
rect 146667 281745 146701 281773
rect 146729 281745 146763 281773
rect 146791 281745 155577 281773
rect 155605 281745 155639 281773
rect 155667 281745 155701 281773
rect 155729 281745 155763 281773
rect 155791 281745 164577 281773
rect 164605 281745 164639 281773
rect 164667 281745 164701 281773
rect 164729 281745 164763 281773
rect 164791 281745 173577 281773
rect 173605 281745 173639 281773
rect 173667 281745 173701 281773
rect 173729 281745 173763 281773
rect 173791 281745 182577 281773
rect 182605 281745 182639 281773
rect 182667 281745 182701 281773
rect 182729 281745 182763 281773
rect 182791 281745 191577 281773
rect 191605 281745 191639 281773
rect 191667 281745 191701 281773
rect 191729 281745 191763 281773
rect 191791 281745 200577 281773
rect 200605 281745 200639 281773
rect 200667 281745 200701 281773
rect 200729 281745 200763 281773
rect 200791 281745 209577 281773
rect 209605 281745 209639 281773
rect 209667 281745 209701 281773
rect 209729 281745 209763 281773
rect 209791 281745 218577 281773
rect 218605 281745 218639 281773
rect 218667 281745 218701 281773
rect 218729 281745 218763 281773
rect 218791 281745 227577 281773
rect 227605 281745 227639 281773
rect 227667 281745 227701 281773
rect 227729 281745 227763 281773
rect 227791 281745 236577 281773
rect 236605 281745 236639 281773
rect 236667 281745 236701 281773
rect 236729 281745 236763 281773
rect 236791 281745 245577 281773
rect 245605 281745 245639 281773
rect 245667 281745 245701 281773
rect 245729 281745 245763 281773
rect 245791 281745 254577 281773
rect 254605 281745 254639 281773
rect 254667 281745 254701 281773
rect 254729 281745 254763 281773
rect 254791 281745 263577 281773
rect 263605 281745 263639 281773
rect 263667 281745 263701 281773
rect 263729 281745 263763 281773
rect 263791 281745 272577 281773
rect 272605 281745 272639 281773
rect 272667 281745 272701 281773
rect 272729 281745 272763 281773
rect 272791 281745 281577 281773
rect 281605 281745 281639 281773
rect 281667 281745 281701 281773
rect 281729 281745 281763 281773
rect 281791 281745 290577 281773
rect 290605 281745 290639 281773
rect 290667 281745 290701 281773
rect 290729 281745 290763 281773
rect 290791 281745 299256 281773
rect 299284 281745 299318 281773
rect 299346 281745 299380 281773
rect 299408 281745 299442 281773
rect 299470 281745 299998 281773
rect -6 281697 299998 281745
rect -6 275959 299998 276007
rect -6 275931 42 275959
rect 70 275931 104 275959
rect 132 275931 166 275959
rect 194 275931 228 275959
rect 256 275931 4437 275959
rect 4465 275931 4499 275959
rect 4527 275931 4561 275959
rect 4589 275931 4623 275959
rect 4651 275931 13437 275959
rect 13465 275931 13499 275959
rect 13527 275931 13561 275959
rect 13589 275931 13623 275959
rect 13651 275931 22437 275959
rect 22465 275931 22499 275959
rect 22527 275931 22561 275959
rect 22589 275931 22623 275959
rect 22651 275931 31437 275959
rect 31465 275931 31499 275959
rect 31527 275931 31561 275959
rect 31589 275931 31623 275959
rect 31651 275931 40437 275959
rect 40465 275931 40499 275959
rect 40527 275931 40561 275959
rect 40589 275931 40623 275959
rect 40651 275931 49437 275959
rect 49465 275931 49499 275959
rect 49527 275931 49561 275959
rect 49589 275931 49623 275959
rect 49651 275931 58437 275959
rect 58465 275931 58499 275959
rect 58527 275931 58561 275959
rect 58589 275931 58623 275959
rect 58651 275931 67437 275959
rect 67465 275931 67499 275959
rect 67527 275931 67561 275959
rect 67589 275931 67623 275959
rect 67651 275931 76437 275959
rect 76465 275931 76499 275959
rect 76527 275931 76561 275959
rect 76589 275931 76623 275959
rect 76651 275931 85437 275959
rect 85465 275931 85499 275959
rect 85527 275931 85561 275959
rect 85589 275931 85623 275959
rect 85651 275931 94437 275959
rect 94465 275931 94499 275959
rect 94527 275931 94561 275959
rect 94589 275931 94623 275959
rect 94651 275931 103437 275959
rect 103465 275931 103499 275959
rect 103527 275931 103561 275959
rect 103589 275931 103623 275959
rect 103651 275931 112437 275959
rect 112465 275931 112499 275959
rect 112527 275931 112561 275959
rect 112589 275931 112623 275959
rect 112651 275931 121437 275959
rect 121465 275931 121499 275959
rect 121527 275931 121561 275959
rect 121589 275931 121623 275959
rect 121651 275931 130437 275959
rect 130465 275931 130499 275959
rect 130527 275931 130561 275959
rect 130589 275931 130623 275959
rect 130651 275931 139437 275959
rect 139465 275931 139499 275959
rect 139527 275931 139561 275959
rect 139589 275931 139623 275959
rect 139651 275931 148437 275959
rect 148465 275931 148499 275959
rect 148527 275931 148561 275959
rect 148589 275931 148623 275959
rect 148651 275931 157437 275959
rect 157465 275931 157499 275959
rect 157527 275931 157561 275959
rect 157589 275931 157623 275959
rect 157651 275931 166437 275959
rect 166465 275931 166499 275959
rect 166527 275931 166561 275959
rect 166589 275931 166623 275959
rect 166651 275931 175437 275959
rect 175465 275931 175499 275959
rect 175527 275931 175561 275959
rect 175589 275931 175623 275959
rect 175651 275931 184437 275959
rect 184465 275931 184499 275959
rect 184527 275931 184561 275959
rect 184589 275931 184623 275959
rect 184651 275931 193437 275959
rect 193465 275931 193499 275959
rect 193527 275931 193561 275959
rect 193589 275931 193623 275959
rect 193651 275931 202437 275959
rect 202465 275931 202499 275959
rect 202527 275931 202561 275959
rect 202589 275931 202623 275959
rect 202651 275931 211437 275959
rect 211465 275931 211499 275959
rect 211527 275931 211561 275959
rect 211589 275931 211623 275959
rect 211651 275931 220437 275959
rect 220465 275931 220499 275959
rect 220527 275931 220561 275959
rect 220589 275931 220623 275959
rect 220651 275931 229437 275959
rect 229465 275931 229499 275959
rect 229527 275931 229561 275959
rect 229589 275931 229623 275959
rect 229651 275931 238437 275959
rect 238465 275931 238499 275959
rect 238527 275931 238561 275959
rect 238589 275931 238623 275959
rect 238651 275931 247437 275959
rect 247465 275931 247499 275959
rect 247527 275931 247561 275959
rect 247589 275931 247623 275959
rect 247651 275931 256437 275959
rect 256465 275931 256499 275959
rect 256527 275931 256561 275959
rect 256589 275931 256623 275959
rect 256651 275931 265437 275959
rect 265465 275931 265499 275959
rect 265527 275931 265561 275959
rect 265589 275931 265623 275959
rect 265651 275931 274437 275959
rect 274465 275931 274499 275959
rect 274527 275931 274561 275959
rect 274589 275931 274623 275959
rect 274651 275931 283437 275959
rect 283465 275931 283499 275959
rect 283527 275931 283561 275959
rect 283589 275931 283623 275959
rect 283651 275931 292437 275959
rect 292465 275931 292499 275959
rect 292527 275931 292561 275959
rect 292589 275931 292623 275959
rect 292651 275931 299736 275959
rect 299764 275931 299798 275959
rect 299826 275931 299860 275959
rect 299888 275931 299922 275959
rect 299950 275931 299998 275959
rect -6 275897 299998 275931
rect -6 275869 42 275897
rect 70 275869 104 275897
rect 132 275869 166 275897
rect 194 275869 228 275897
rect 256 275869 4437 275897
rect 4465 275869 4499 275897
rect 4527 275869 4561 275897
rect 4589 275869 4623 275897
rect 4651 275869 13437 275897
rect 13465 275869 13499 275897
rect 13527 275869 13561 275897
rect 13589 275869 13623 275897
rect 13651 275869 22437 275897
rect 22465 275869 22499 275897
rect 22527 275869 22561 275897
rect 22589 275869 22623 275897
rect 22651 275869 31437 275897
rect 31465 275869 31499 275897
rect 31527 275869 31561 275897
rect 31589 275869 31623 275897
rect 31651 275869 40437 275897
rect 40465 275869 40499 275897
rect 40527 275869 40561 275897
rect 40589 275869 40623 275897
rect 40651 275869 49437 275897
rect 49465 275869 49499 275897
rect 49527 275869 49561 275897
rect 49589 275869 49623 275897
rect 49651 275869 58437 275897
rect 58465 275869 58499 275897
rect 58527 275869 58561 275897
rect 58589 275869 58623 275897
rect 58651 275869 67437 275897
rect 67465 275869 67499 275897
rect 67527 275869 67561 275897
rect 67589 275869 67623 275897
rect 67651 275869 76437 275897
rect 76465 275869 76499 275897
rect 76527 275869 76561 275897
rect 76589 275869 76623 275897
rect 76651 275869 85437 275897
rect 85465 275869 85499 275897
rect 85527 275869 85561 275897
rect 85589 275869 85623 275897
rect 85651 275869 94437 275897
rect 94465 275869 94499 275897
rect 94527 275869 94561 275897
rect 94589 275869 94623 275897
rect 94651 275869 103437 275897
rect 103465 275869 103499 275897
rect 103527 275869 103561 275897
rect 103589 275869 103623 275897
rect 103651 275869 112437 275897
rect 112465 275869 112499 275897
rect 112527 275869 112561 275897
rect 112589 275869 112623 275897
rect 112651 275869 121437 275897
rect 121465 275869 121499 275897
rect 121527 275869 121561 275897
rect 121589 275869 121623 275897
rect 121651 275869 130437 275897
rect 130465 275869 130499 275897
rect 130527 275869 130561 275897
rect 130589 275869 130623 275897
rect 130651 275869 139437 275897
rect 139465 275869 139499 275897
rect 139527 275869 139561 275897
rect 139589 275869 139623 275897
rect 139651 275869 148437 275897
rect 148465 275869 148499 275897
rect 148527 275869 148561 275897
rect 148589 275869 148623 275897
rect 148651 275869 157437 275897
rect 157465 275869 157499 275897
rect 157527 275869 157561 275897
rect 157589 275869 157623 275897
rect 157651 275869 166437 275897
rect 166465 275869 166499 275897
rect 166527 275869 166561 275897
rect 166589 275869 166623 275897
rect 166651 275869 175437 275897
rect 175465 275869 175499 275897
rect 175527 275869 175561 275897
rect 175589 275869 175623 275897
rect 175651 275869 184437 275897
rect 184465 275869 184499 275897
rect 184527 275869 184561 275897
rect 184589 275869 184623 275897
rect 184651 275869 193437 275897
rect 193465 275869 193499 275897
rect 193527 275869 193561 275897
rect 193589 275869 193623 275897
rect 193651 275869 202437 275897
rect 202465 275869 202499 275897
rect 202527 275869 202561 275897
rect 202589 275869 202623 275897
rect 202651 275869 211437 275897
rect 211465 275869 211499 275897
rect 211527 275869 211561 275897
rect 211589 275869 211623 275897
rect 211651 275869 220437 275897
rect 220465 275869 220499 275897
rect 220527 275869 220561 275897
rect 220589 275869 220623 275897
rect 220651 275869 229437 275897
rect 229465 275869 229499 275897
rect 229527 275869 229561 275897
rect 229589 275869 229623 275897
rect 229651 275869 238437 275897
rect 238465 275869 238499 275897
rect 238527 275869 238561 275897
rect 238589 275869 238623 275897
rect 238651 275869 247437 275897
rect 247465 275869 247499 275897
rect 247527 275869 247561 275897
rect 247589 275869 247623 275897
rect 247651 275869 256437 275897
rect 256465 275869 256499 275897
rect 256527 275869 256561 275897
rect 256589 275869 256623 275897
rect 256651 275869 265437 275897
rect 265465 275869 265499 275897
rect 265527 275869 265561 275897
rect 265589 275869 265623 275897
rect 265651 275869 274437 275897
rect 274465 275869 274499 275897
rect 274527 275869 274561 275897
rect 274589 275869 274623 275897
rect 274651 275869 283437 275897
rect 283465 275869 283499 275897
rect 283527 275869 283561 275897
rect 283589 275869 283623 275897
rect 283651 275869 292437 275897
rect 292465 275869 292499 275897
rect 292527 275869 292561 275897
rect 292589 275869 292623 275897
rect 292651 275869 299736 275897
rect 299764 275869 299798 275897
rect 299826 275869 299860 275897
rect 299888 275869 299922 275897
rect 299950 275869 299998 275897
rect -6 275835 299998 275869
rect -6 275807 42 275835
rect 70 275807 104 275835
rect 132 275807 166 275835
rect 194 275807 228 275835
rect 256 275807 4437 275835
rect 4465 275807 4499 275835
rect 4527 275807 4561 275835
rect 4589 275807 4623 275835
rect 4651 275807 13437 275835
rect 13465 275807 13499 275835
rect 13527 275807 13561 275835
rect 13589 275807 13623 275835
rect 13651 275807 22437 275835
rect 22465 275807 22499 275835
rect 22527 275807 22561 275835
rect 22589 275807 22623 275835
rect 22651 275807 31437 275835
rect 31465 275807 31499 275835
rect 31527 275807 31561 275835
rect 31589 275807 31623 275835
rect 31651 275807 40437 275835
rect 40465 275807 40499 275835
rect 40527 275807 40561 275835
rect 40589 275807 40623 275835
rect 40651 275807 49437 275835
rect 49465 275807 49499 275835
rect 49527 275807 49561 275835
rect 49589 275807 49623 275835
rect 49651 275807 58437 275835
rect 58465 275807 58499 275835
rect 58527 275807 58561 275835
rect 58589 275807 58623 275835
rect 58651 275807 67437 275835
rect 67465 275807 67499 275835
rect 67527 275807 67561 275835
rect 67589 275807 67623 275835
rect 67651 275807 76437 275835
rect 76465 275807 76499 275835
rect 76527 275807 76561 275835
rect 76589 275807 76623 275835
rect 76651 275807 85437 275835
rect 85465 275807 85499 275835
rect 85527 275807 85561 275835
rect 85589 275807 85623 275835
rect 85651 275807 94437 275835
rect 94465 275807 94499 275835
rect 94527 275807 94561 275835
rect 94589 275807 94623 275835
rect 94651 275807 103437 275835
rect 103465 275807 103499 275835
rect 103527 275807 103561 275835
rect 103589 275807 103623 275835
rect 103651 275807 112437 275835
rect 112465 275807 112499 275835
rect 112527 275807 112561 275835
rect 112589 275807 112623 275835
rect 112651 275807 121437 275835
rect 121465 275807 121499 275835
rect 121527 275807 121561 275835
rect 121589 275807 121623 275835
rect 121651 275807 130437 275835
rect 130465 275807 130499 275835
rect 130527 275807 130561 275835
rect 130589 275807 130623 275835
rect 130651 275807 139437 275835
rect 139465 275807 139499 275835
rect 139527 275807 139561 275835
rect 139589 275807 139623 275835
rect 139651 275807 148437 275835
rect 148465 275807 148499 275835
rect 148527 275807 148561 275835
rect 148589 275807 148623 275835
rect 148651 275807 157437 275835
rect 157465 275807 157499 275835
rect 157527 275807 157561 275835
rect 157589 275807 157623 275835
rect 157651 275807 166437 275835
rect 166465 275807 166499 275835
rect 166527 275807 166561 275835
rect 166589 275807 166623 275835
rect 166651 275807 175437 275835
rect 175465 275807 175499 275835
rect 175527 275807 175561 275835
rect 175589 275807 175623 275835
rect 175651 275807 184437 275835
rect 184465 275807 184499 275835
rect 184527 275807 184561 275835
rect 184589 275807 184623 275835
rect 184651 275807 193437 275835
rect 193465 275807 193499 275835
rect 193527 275807 193561 275835
rect 193589 275807 193623 275835
rect 193651 275807 202437 275835
rect 202465 275807 202499 275835
rect 202527 275807 202561 275835
rect 202589 275807 202623 275835
rect 202651 275807 211437 275835
rect 211465 275807 211499 275835
rect 211527 275807 211561 275835
rect 211589 275807 211623 275835
rect 211651 275807 220437 275835
rect 220465 275807 220499 275835
rect 220527 275807 220561 275835
rect 220589 275807 220623 275835
rect 220651 275807 229437 275835
rect 229465 275807 229499 275835
rect 229527 275807 229561 275835
rect 229589 275807 229623 275835
rect 229651 275807 238437 275835
rect 238465 275807 238499 275835
rect 238527 275807 238561 275835
rect 238589 275807 238623 275835
rect 238651 275807 247437 275835
rect 247465 275807 247499 275835
rect 247527 275807 247561 275835
rect 247589 275807 247623 275835
rect 247651 275807 256437 275835
rect 256465 275807 256499 275835
rect 256527 275807 256561 275835
rect 256589 275807 256623 275835
rect 256651 275807 265437 275835
rect 265465 275807 265499 275835
rect 265527 275807 265561 275835
rect 265589 275807 265623 275835
rect 265651 275807 274437 275835
rect 274465 275807 274499 275835
rect 274527 275807 274561 275835
rect 274589 275807 274623 275835
rect 274651 275807 283437 275835
rect 283465 275807 283499 275835
rect 283527 275807 283561 275835
rect 283589 275807 283623 275835
rect 283651 275807 292437 275835
rect 292465 275807 292499 275835
rect 292527 275807 292561 275835
rect 292589 275807 292623 275835
rect 292651 275807 299736 275835
rect 299764 275807 299798 275835
rect 299826 275807 299860 275835
rect 299888 275807 299922 275835
rect 299950 275807 299998 275835
rect -6 275773 299998 275807
rect -6 275745 42 275773
rect 70 275745 104 275773
rect 132 275745 166 275773
rect 194 275745 228 275773
rect 256 275745 4437 275773
rect 4465 275745 4499 275773
rect 4527 275745 4561 275773
rect 4589 275745 4623 275773
rect 4651 275745 13437 275773
rect 13465 275745 13499 275773
rect 13527 275745 13561 275773
rect 13589 275745 13623 275773
rect 13651 275745 22437 275773
rect 22465 275745 22499 275773
rect 22527 275745 22561 275773
rect 22589 275745 22623 275773
rect 22651 275745 31437 275773
rect 31465 275745 31499 275773
rect 31527 275745 31561 275773
rect 31589 275745 31623 275773
rect 31651 275745 40437 275773
rect 40465 275745 40499 275773
rect 40527 275745 40561 275773
rect 40589 275745 40623 275773
rect 40651 275745 49437 275773
rect 49465 275745 49499 275773
rect 49527 275745 49561 275773
rect 49589 275745 49623 275773
rect 49651 275745 58437 275773
rect 58465 275745 58499 275773
rect 58527 275745 58561 275773
rect 58589 275745 58623 275773
rect 58651 275745 67437 275773
rect 67465 275745 67499 275773
rect 67527 275745 67561 275773
rect 67589 275745 67623 275773
rect 67651 275745 76437 275773
rect 76465 275745 76499 275773
rect 76527 275745 76561 275773
rect 76589 275745 76623 275773
rect 76651 275745 85437 275773
rect 85465 275745 85499 275773
rect 85527 275745 85561 275773
rect 85589 275745 85623 275773
rect 85651 275745 94437 275773
rect 94465 275745 94499 275773
rect 94527 275745 94561 275773
rect 94589 275745 94623 275773
rect 94651 275745 103437 275773
rect 103465 275745 103499 275773
rect 103527 275745 103561 275773
rect 103589 275745 103623 275773
rect 103651 275745 112437 275773
rect 112465 275745 112499 275773
rect 112527 275745 112561 275773
rect 112589 275745 112623 275773
rect 112651 275745 121437 275773
rect 121465 275745 121499 275773
rect 121527 275745 121561 275773
rect 121589 275745 121623 275773
rect 121651 275745 130437 275773
rect 130465 275745 130499 275773
rect 130527 275745 130561 275773
rect 130589 275745 130623 275773
rect 130651 275745 139437 275773
rect 139465 275745 139499 275773
rect 139527 275745 139561 275773
rect 139589 275745 139623 275773
rect 139651 275745 148437 275773
rect 148465 275745 148499 275773
rect 148527 275745 148561 275773
rect 148589 275745 148623 275773
rect 148651 275745 157437 275773
rect 157465 275745 157499 275773
rect 157527 275745 157561 275773
rect 157589 275745 157623 275773
rect 157651 275745 166437 275773
rect 166465 275745 166499 275773
rect 166527 275745 166561 275773
rect 166589 275745 166623 275773
rect 166651 275745 175437 275773
rect 175465 275745 175499 275773
rect 175527 275745 175561 275773
rect 175589 275745 175623 275773
rect 175651 275745 184437 275773
rect 184465 275745 184499 275773
rect 184527 275745 184561 275773
rect 184589 275745 184623 275773
rect 184651 275745 193437 275773
rect 193465 275745 193499 275773
rect 193527 275745 193561 275773
rect 193589 275745 193623 275773
rect 193651 275745 202437 275773
rect 202465 275745 202499 275773
rect 202527 275745 202561 275773
rect 202589 275745 202623 275773
rect 202651 275745 211437 275773
rect 211465 275745 211499 275773
rect 211527 275745 211561 275773
rect 211589 275745 211623 275773
rect 211651 275745 220437 275773
rect 220465 275745 220499 275773
rect 220527 275745 220561 275773
rect 220589 275745 220623 275773
rect 220651 275745 229437 275773
rect 229465 275745 229499 275773
rect 229527 275745 229561 275773
rect 229589 275745 229623 275773
rect 229651 275745 238437 275773
rect 238465 275745 238499 275773
rect 238527 275745 238561 275773
rect 238589 275745 238623 275773
rect 238651 275745 247437 275773
rect 247465 275745 247499 275773
rect 247527 275745 247561 275773
rect 247589 275745 247623 275773
rect 247651 275745 256437 275773
rect 256465 275745 256499 275773
rect 256527 275745 256561 275773
rect 256589 275745 256623 275773
rect 256651 275745 265437 275773
rect 265465 275745 265499 275773
rect 265527 275745 265561 275773
rect 265589 275745 265623 275773
rect 265651 275745 274437 275773
rect 274465 275745 274499 275773
rect 274527 275745 274561 275773
rect 274589 275745 274623 275773
rect 274651 275745 283437 275773
rect 283465 275745 283499 275773
rect 283527 275745 283561 275773
rect 283589 275745 283623 275773
rect 283651 275745 292437 275773
rect 292465 275745 292499 275773
rect 292527 275745 292561 275773
rect 292589 275745 292623 275773
rect 292651 275745 299736 275773
rect 299764 275745 299798 275773
rect 299826 275745 299860 275773
rect 299888 275745 299922 275773
rect 299950 275745 299998 275773
rect -6 275697 299998 275745
rect -6 272959 299998 273007
rect -6 272931 522 272959
rect 550 272931 584 272959
rect 612 272931 646 272959
rect 674 272931 708 272959
rect 736 272931 2577 272959
rect 2605 272931 2639 272959
rect 2667 272931 2701 272959
rect 2729 272931 2763 272959
rect 2791 272931 11577 272959
rect 11605 272931 11639 272959
rect 11667 272931 11701 272959
rect 11729 272931 11763 272959
rect 11791 272931 20577 272959
rect 20605 272931 20639 272959
rect 20667 272931 20701 272959
rect 20729 272931 20763 272959
rect 20791 272931 29577 272959
rect 29605 272931 29639 272959
rect 29667 272931 29701 272959
rect 29729 272931 29763 272959
rect 29791 272931 38577 272959
rect 38605 272931 38639 272959
rect 38667 272931 38701 272959
rect 38729 272931 38763 272959
rect 38791 272931 47577 272959
rect 47605 272931 47639 272959
rect 47667 272931 47701 272959
rect 47729 272931 47763 272959
rect 47791 272931 56577 272959
rect 56605 272931 56639 272959
rect 56667 272931 56701 272959
rect 56729 272931 56763 272959
rect 56791 272931 65577 272959
rect 65605 272931 65639 272959
rect 65667 272931 65701 272959
rect 65729 272931 65763 272959
rect 65791 272931 74577 272959
rect 74605 272931 74639 272959
rect 74667 272931 74701 272959
rect 74729 272931 74763 272959
rect 74791 272931 83577 272959
rect 83605 272931 83639 272959
rect 83667 272931 83701 272959
rect 83729 272931 83763 272959
rect 83791 272931 92577 272959
rect 92605 272931 92639 272959
rect 92667 272931 92701 272959
rect 92729 272931 92763 272959
rect 92791 272931 101577 272959
rect 101605 272931 101639 272959
rect 101667 272931 101701 272959
rect 101729 272931 101763 272959
rect 101791 272931 110577 272959
rect 110605 272931 110639 272959
rect 110667 272931 110701 272959
rect 110729 272931 110763 272959
rect 110791 272931 119577 272959
rect 119605 272931 119639 272959
rect 119667 272931 119701 272959
rect 119729 272931 119763 272959
rect 119791 272931 128577 272959
rect 128605 272931 128639 272959
rect 128667 272931 128701 272959
rect 128729 272931 128763 272959
rect 128791 272931 137577 272959
rect 137605 272931 137639 272959
rect 137667 272931 137701 272959
rect 137729 272931 137763 272959
rect 137791 272931 146577 272959
rect 146605 272931 146639 272959
rect 146667 272931 146701 272959
rect 146729 272931 146763 272959
rect 146791 272931 155577 272959
rect 155605 272931 155639 272959
rect 155667 272931 155701 272959
rect 155729 272931 155763 272959
rect 155791 272931 164577 272959
rect 164605 272931 164639 272959
rect 164667 272931 164701 272959
rect 164729 272931 164763 272959
rect 164791 272931 173577 272959
rect 173605 272931 173639 272959
rect 173667 272931 173701 272959
rect 173729 272931 173763 272959
rect 173791 272931 182577 272959
rect 182605 272931 182639 272959
rect 182667 272931 182701 272959
rect 182729 272931 182763 272959
rect 182791 272931 191577 272959
rect 191605 272931 191639 272959
rect 191667 272931 191701 272959
rect 191729 272931 191763 272959
rect 191791 272931 200577 272959
rect 200605 272931 200639 272959
rect 200667 272931 200701 272959
rect 200729 272931 200763 272959
rect 200791 272931 209577 272959
rect 209605 272931 209639 272959
rect 209667 272931 209701 272959
rect 209729 272931 209763 272959
rect 209791 272931 218577 272959
rect 218605 272931 218639 272959
rect 218667 272931 218701 272959
rect 218729 272931 218763 272959
rect 218791 272931 227577 272959
rect 227605 272931 227639 272959
rect 227667 272931 227701 272959
rect 227729 272931 227763 272959
rect 227791 272931 236577 272959
rect 236605 272931 236639 272959
rect 236667 272931 236701 272959
rect 236729 272931 236763 272959
rect 236791 272931 245577 272959
rect 245605 272931 245639 272959
rect 245667 272931 245701 272959
rect 245729 272931 245763 272959
rect 245791 272931 254577 272959
rect 254605 272931 254639 272959
rect 254667 272931 254701 272959
rect 254729 272931 254763 272959
rect 254791 272931 263577 272959
rect 263605 272931 263639 272959
rect 263667 272931 263701 272959
rect 263729 272931 263763 272959
rect 263791 272931 272577 272959
rect 272605 272931 272639 272959
rect 272667 272931 272701 272959
rect 272729 272931 272763 272959
rect 272791 272931 281577 272959
rect 281605 272931 281639 272959
rect 281667 272931 281701 272959
rect 281729 272931 281763 272959
rect 281791 272931 290577 272959
rect 290605 272931 290639 272959
rect 290667 272931 290701 272959
rect 290729 272931 290763 272959
rect 290791 272931 299256 272959
rect 299284 272931 299318 272959
rect 299346 272931 299380 272959
rect 299408 272931 299442 272959
rect 299470 272931 299998 272959
rect -6 272897 299998 272931
rect -6 272869 522 272897
rect 550 272869 584 272897
rect 612 272869 646 272897
rect 674 272869 708 272897
rect 736 272869 2577 272897
rect 2605 272869 2639 272897
rect 2667 272869 2701 272897
rect 2729 272869 2763 272897
rect 2791 272869 11577 272897
rect 11605 272869 11639 272897
rect 11667 272869 11701 272897
rect 11729 272869 11763 272897
rect 11791 272869 20577 272897
rect 20605 272869 20639 272897
rect 20667 272869 20701 272897
rect 20729 272869 20763 272897
rect 20791 272869 29577 272897
rect 29605 272869 29639 272897
rect 29667 272869 29701 272897
rect 29729 272869 29763 272897
rect 29791 272869 38577 272897
rect 38605 272869 38639 272897
rect 38667 272869 38701 272897
rect 38729 272869 38763 272897
rect 38791 272869 47577 272897
rect 47605 272869 47639 272897
rect 47667 272869 47701 272897
rect 47729 272869 47763 272897
rect 47791 272869 56577 272897
rect 56605 272869 56639 272897
rect 56667 272869 56701 272897
rect 56729 272869 56763 272897
rect 56791 272869 65577 272897
rect 65605 272869 65639 272897
rect 65667 272869 65701 272897
rect 65729 272869 65763 272897
rect 65791 272869 74577 272897
rect 74605 272869 74639 272897
rect 74667 272869 74701 272897
rect 74729 272869 74763 272897
rect 74791 272869 83577 272897
rect 83605 272869 83639 272897
rect 83667 272869 83701 272897
rect 83729 272869 83763 272897
rect 83791 272869 92577 272897
rect 92605 272869 92639 272897
rect 92667 272869 92701 272897
rect 92729 272869 92763 272897
rect 92791 272869 101577 272897
rect 101605 272869 101639 272897
rect 101667 272869 101701 272897
rect 101729 272869 101763 272897
rect 101791 272869 110577 272897
rect 110605 272869 110639 272897
rect 110667 272869 110701 272897
rect 110729 272869 110763 272897
rect 110791 272869 119577 272897
rect 119605 272869 119639 272897
rect 119667 272869 119701 272897
rect 119729 272869 119763 272897
rect 119791 272869 128577 272897
rect 128605 272869 128639 272897
rect 128667 272869 128701 272897
rect 128729 272869 128763 272897
rect 128791 272869 137577 272897
rect 137605 272869 137639 272897
rect 137667 272869 137701 272897
rect 137729 272869 137763 272897
rect 137791 272869 146577 272897
rect 146605 272869 146639 272897
rect 146667 272869 146701 272897
rect 146729 272869 146763 272897
rect 146791 272869 155577 272897
rect 155605 272869 155639 272897
rect 155667 272869 155701 272897
rect 155729 272869 155763 272897
rect 155791 272869 164577 272897
rect 164605 272869 164639 272897
rect 164667 272869 164701 272897
rect 164729 272869 164763 272897
rect 164791 272869 173577 272897
rect 173605 272869 173639 272897
rect 173667 272869 173701 272897
rect 173729 272869 173763 272897
rect 173791 272869 182577 272897
rect 182605 272869 182639 272897
rect 182667 272869 182701 272897
rect 182729 272869 182763 272897
rect 182791 272869 191577 272897
rect 191605 272869 191639 272897
rect 191667 272869 191701 272897
rect 191729 272869 191763 272897
rect 191791 272869 200577 272897
rect 200605 272869 200639 272897
rect 200667 272869 200701 272897
rect 200729 272869 200763 272897
rect 200791 272869 209577 272897
rect 209605 272869 209639 272897
rect 209667 272869 209701 272897
rect 209729 272869 209763 272897
rect 209791 272869 218577 272897
rect 218605 272869 218639 272897
rect 218667 272869 218701 272897
rect 218729 272869 218763 272897
rect 218791 272869 227577 272897
rect 227605 272869 227639 272897
rect 227667 272869 227701 272897
rect 227729 272869 227763 272897
rect 227791 272869 236577 272897
rect 236605 272869 236639 272897
rect 236667 272869 236701 272897
rect 236729 272869 236763 272897
rect 236791 272869 245577 272897
rect 245605 272869 245639 272897
rect 245667 272869 245701 272897
rect 245729 272869 245763 272897
rect 245791 272869 254577 272897
rect 254605 272869 254639 272897
rect 254667 272869 254701 272897
rect 254729 272869 254763 272897
rect 254791 272869 263577 272897
rect 263605 272869 263639 272897
rect 263667 272869 263701 272897
rect 263729 272869 263763 272897
rect 263791 272869 272577 272897
rect 272605 272869 272639 272897
rect 272667 272869 272701 272897
rect 272729 272869 272763 272897
rect 272791 272869 281577 272897
rect 281605 272869 281639 272897
rect 281667 272869 281701 272897
rect 281729 272869 281763 272897
rect 281791 272869 290577 272897
rect 290605 272869 290639 272897
rect 290667 272869 290701 272897
rect 290729 272869 290763 272897
rect 290791 272869 299256 272897
rect 299284 272869 299318 272897
rect 299346 272869 299380 272897
rect 299408 272869 299442 272897
rect 299470 272869 299998 272897
rect -6 272835 299998 272869
rect -6 272807 522 272835
rect 550 272807 584 272835
rect 612 272807 646 272835
rect 674 272807 708 272835
rect 736 272807 2577 272835
rect 2605 272807 2639 272835
rect 2667 272807 2701 272835
rect 2729 272807 2763 272835
rect 2791 272807 11577 272835
rect 11605 272807 11639 272835
rect 11667 272807 11701 272835
rect 11729 272807 11763 272835
rect 11791 272807 20577 272835
rect 20605 272807 20639 272835
rect 20667 272807 20701 272835
rect 20729 272807 20763 272835
rect 20791 272807 29577 272835
rect 29605 272807 29639 272835
rect 29667 272807 29701 272835
rect 29729 272807 29763 272835
rect 29791 272807 38577 272835
rect 38605 272807 38639 272835
rect 38667 272807 38701 272835
rect 38729 272807 38763 272835
rect 38791 272807 47577 272835
rect 47605 272807 47639 272835
rect 47667 272807 47701 272835
rect 47729 272807 47763 272835
rect 47791 272807 56577 272835
rect 56605 272807 56639 272835
rect 56667 272807 56701 272835
rect 56729 272807 56763 272835
rect 56791 272807 65577 272835
rect 65605 272807 65639 272835
rect 65667 272807 65701 272835
rect 65729 272807 65763 272835
rect 65791 272807 74577 272835
rect 74605 272807 74639 272835
rect 74667 272807 74701 272835
rect 74729 272807 74763 272835
rect 74791 272807 83577 272835
rect 83605 272807 83639 272835
rect 83667 272807 83701 272835
rect 83729 272807 83763 272835
rect 83791 272807 92577 272835
rect 92605 272807 92639 272835
rect 92667 272807 92701 272835
rect 92729 272807 92763 272835
rect 92791 272807 101577 272835
rect 101605 272807 101639 272835
rect 101667 272807 101701 272835
rect 101729 272807 101763 272835
rect 101791 272807 110577 272835
rect 110605 272807 110639 272835
rect 110667 272807 110701 272835
rect 110729 272807 110763 272835
rect 110791 272807 119577 272835
rect 119605 272807 119639 272835
rect 119667 272807 119701 272835
rect 119729 272807 119763 272835
rect 119791 272807 128577 272835
rect 128605 272807 128639 272835
rect 128667 272807 128701 272835
rect 128729 272807 128763 272835
rect 128791 272807 137577 272835
rect 137605 272807 137639 272835
rect 137667 272807 137701 272835
rect 137729 272807 137763 272835
rect 137791 272807 146577 272835
rect 146605 272807 146639 272835
rect 146667 272807 146701 272835
rect 146729 272807 146763 272835
rect 146791 272807 155577 272835
rect 155605 272807 155639 272835
rect 155667 272807 155701 272835
rect 155729 272807 155763 272835
rect 155791 272807 164577 272835
rect 164605 272807 164639 272835
rect 164667 272807 164701 272835
rect 164729 272807 164763 272835
rect 164791 272807 173577 272835
rect 173605 272807 173639 272835
rect 173667 272807 173701 272835
rect 173729 272807 173763 272835
rect 173791 272807 182577 272835
rect 182605 272807 182639 272835
rect 182667 272807 182701 272835
rect 182729 272807 182763 272835
rect 182791 272807 191577 272835
rect 191605 272807 191639 272835
rect 191667 272807 191701 272835
rect 191729 272807 191763 272835
rect 191791 272807 200577 272835
rect 200605 272807 200639 272835
rect 200667 272807 200701 272835
rect 200729 272807 200763 272835
rect 200791 272807 209577 272835
rect 209605 272807 209639 272835
rect 209667 272807 209701 272835
rect 209729 272807 209763 272835
rect 209791 272807 218577 272835
rect 218605 272807 218639 272835
rect 218667 272807 218701 272835
rect 218729 272807 218763 272835
rect 218791 272807 227577 272835
rect 227605 272807 227639 272835
rect 227667 272807 227701 272835
rect 227729 272807 227763 272835
rect 227791 272807 236577 272835
rect 236605 272807 236639 272835
rect 236667 272807 236701 272835
rect 236729 272807 236763 272835
rect 236791 272807 245577 272835
rect 245605 272807 245639 272835
rect 245667 272807 245701 272835
rect 245729 272807 245763 272835
rect 245791 272807 254577 272835
rect 254605 272807 254639 272835
rect 254667 272807 254701 272835
rect 254729 272807 254763 272835
rect 254791 272807 263577 272835
rect 263605 272807 263639 272835
rect 263667 272807 263701 272835
rect 263729 272807 263763 272835
rect 263791 272807 272577 272835
rect 272605 272807 272639 272835
rect 272667 272807 272701 272835
rect 272729 272807 272763 272835
rect 272791 272807 281577 272835
rect 281605 272807 281639 272835
rect 281667 272807 281701 272835
rect 281729 272807 281763 272835
rect 281791 272807 290577 272835
rect 290605 272807 290639 272835
rect 290667 272807 290701 272835
rect 290729 272807 290763 272835
rect 290791 272807 299256 272835
rect 299284 272807 299318 272835
rect 299346 272807 299380 272835
rect 299408 272807 299442 272835
rect 299470 272807 299998 272835
rect -6 272773 299998 272807
rect -6 272745 522 272773
rect 550 272745 584 272773
rect 612 272745 646 272773
rect 674 272745 708 272773
rect 736 272745 2577 272773
rect 2605 272745 2639 272773
rect 2667 272745 2701 272773
rect 2729 272745 2763 272773
rect 2791 272745 11577 272773
rect 11605 272745 11639 272773
rect 11667 272745 11701 272773
rect 11729 272745 11763 272773
rect 11791 272745 20577 272773
rect 20605 272745 20639 272773
rect 20667 272745 20701 272773
rect 20729 272745 20763 272773
rect 20791 272745 29577 272773
rect 29605 272745 29639 272773
rect 29667 272745 29701 272773
rect 29729 272745 29763 272773
rect 29791 272745 38577 272773
rect 38605 272745 38639 272773
rect 38667 272745 38701 272773
rect 38729 272745 38763 272773
rect 38791 272745 47577 272773
rect 47605 272745 47639 272773
rect 47667 272745 47701 272773
rect 47729 272745 47763 272773
rect 47791 272745 56577 272773
rect 56605 272745 56639 272773
rect 56667 272745 56701 272773
rect 56729 272745 56763 272773
rect 56791 272745 65577 272773
rect 65605 272745 65639 272773
rect 65667 272745 65701 272773
rect 65729 272745 65763 272773
rect 65791 272745 74577 272773
rect 74605 272745 74639 272773
rect 74667 272745 74701 272773
rect 74729 272745 74763 272773
rect 74791 272745 83577 272773
rect 83605 272745 83639 272773
rect 83667 272745 83701 272773
rect 83729 272745 83763 272773
rect 83791 272745 92577 272773
rect 92605 272745 92639 272773
rect 92667 272745 92701 272773
rect 92729 272745 92763 272773
rect 92791 272745 101577 272773
rect 101605 272745 101639 272773
rect 101667 272745 101701 272773
rect 101729 272745 101763 272773
rect 101791 272745 110577 272773
rect 110605 272745 110639 272773
rect 110667 272745 110701 272773
rect 110729 272745 110763 272773
rect 110791 272745 119577 272773
rect 119605 272745 119639 272773
rect 119667 272745 119701 272773
rect 119729 272745 119763 272773
rect 119791 272745 128577 272773
rect 128605 272745 128639 272773
rect 128667 272745 128701 272773
rect 128729 272745 128763 272773
rect 128791 272745 137577 272773
rect 137605 272745 137639 272773
rect 137667 272745 137701 272773
rect 137729 272745 137763 272773
rect 137791 272745 146577 272773
rect 146605 272745 146639 272773
rect 146667 272745 146701 272773
rect 146729 272745 146763 272773
rect 146791 272745 155577 272773
rect 155605 272745 155639 272773
rect 155667 272745 155701 272773
rect 155729 272745 155763 272773
rect 155791 272745 164577 272773
rect 164605 272745 164639 272773
rect 164667 272745 164701 272773
rect 164729 272745 164763 272773
rect 164791 272745 173577 272773
rect 173605 272745 173639 272773
rect 173667 272745 173701 272773
rect 173729 272745 173763 272773
rect 173791 272745 182577 272773
rect 182605 272745 182639 272773
rect 182667 272745 182701 272773
rect 182729 272745 182763 272773
rect 182791 272745 191577 272773
rect 191605 272745 191639 272773
rect 191667 272745 191701 272773
rect 191729 272745 191763 272773
rect 191791 272745 200577 272773
rect 200605 272745 200639 272773
rect 200667 272745 200701 272773
rect 200729 272745 200763 272773
rect 200791 272745 209577 272773
rect 209605 272745 209639 272773
rect 209667 272745 209701 272773
rect 209729 272745 209763 272773
rect 209791 272745 218577 272773
rect 218605 272745 218639 272773
rect 218667 272745 218701 272773
rect 218729 272745 218763 272773
rect 218791 272745 227577 272773
rect 227605 272745 227639 272773
rect 227667 272745 227701 272773
rect 227729 272745 227763 272773
rect 227791 272745 236577 272773
rect 236605 272745 236639 272773
rect 236667 272745 236701 272773
rect 236729 272745 236763 272773
rect 236791 272745 245577 272773
rect 245605 272745 245639 272773
rect 245667 272745 245701 272773
rect 245729 272745 245763 272773
rect 245791 272745 254577 272773
rect 254605 272745 254639 272773
rect 254667 272745 254701 272773
rect 254729 272745 254763 272773
rect 254791 272745 263577 272773
rect 263605 272745 263639 272773
rect 263667 272745 263701 272773
rect 263729 272745 263763 272773
rect 263791 272745 272577 272773
rect 272605 272745 272639 272773
rect 272667 272745 272701 272773
rect 272729 272745 272763 272773
rect 272791 272745 281577 272773
rect 281605 272745 281639 272773
rect 281667 272745 281701 272773
rect 281729 272745 281763 272773
rect 281791 272745 290577 272773
rect 290605 272745 290639 272773
rect 290667 272745 290701 272773
rect 290729 272745 290763 272773
rect 290791 272745 299256 272773
rect 299284 272745 299318 272773
rect 299346 272745 299380 272773
rect 299408 272745 299442 272773
rect 299470 272745 299998 272773
rect -6 272697 299998 272745
rect -6 266959 299998 267007
rect -6 266931 42 266959
rect 70 266931 104 266959
rect 132 266931 166 266959
rect 194 266931 228 266959
rect 256 266931 4437 266959
rect 4465 266931 4499 266959
rect 4527 266931 4561 266959
rect 4589 266931 4623 266959
rect 4651 266931 13437 266959
rect 13465 266931 13499 266959
rect 13527 266931 13561 266959
rect 13589 266931 13623 266959
rect 13651 266931 22437 266959
rect 22465 266931 22499 266959
rect 22527 266931 22561 266959
rect 22589 266931 22623 266959
rect 22651 266931 31437 266959
rect 31465 266931 31499 266959
rect 31527 266931 31561 266959
rect 31589 266931 31623 266959
rect 31651 266931 40437 266959
rect 40465 266931 40499 266959
rect 40527 266931 40561 266959
rect 40589 266931 40623 266959
rect 40651 266931 49437 266959
rect 49465 266931 49499 266959
rect 49527 266931 49561 266959
rect 49589 266931 49623 266959
rect 49651 266931 58437 266959
rect 58465 266931 58499 266959
rect 58527 266931 58561 266959
rect 58589 266931 58623 266959
rect 58651 266931 67437 266959
rect 67465 266931 67499 266959
rect 67527 266931 67561 266959
rect 67589 266931 67623 266959
rect 67651 266931 76437 266959
rect 76465 266931 76499 266959
rect 76527 266931 76561 266959
rect 76589 266931 76623 266959
rect 76651 266931 85437 266959
rect 85465 266931 85499 266959
rect 85527 266931 85561 266959
rect 85589 266931 85623 266959
rect 85651 266931 94437 266959
rect 94465 266931 94499 266959
rect 94527 266931 94561 266959
rect 94589 266931 94623 266959
rect 94651 266931 103437 266959
rect 103465 266931 103499 266959
rect 103527 266931 103561 266959
rect 103589 266931 103623 266959
rect 103651 266931 112437 266959
rect 112465 266931 112499 266959
rect 112527 266931 112561 266959
rect 112589 266931 112623 266959
rect 112651 266931 121437 266959
rect 121465 266931 121499 266959
rect 121527 266931 121561 266959
rect 121589 266931 121623 266959
rect 121651 266931 130437 266959
rect 130465 266931 130499 266959
rect 130527 266931 130561 266959
rect 130589 266931 130623 266959
rect 130651 266931 139437 266959
rect 139465 266931 139499 266959
rect 139527 266931 139561 266959
rect 139589 266931 139623 266959
rect 139651 266931 148437 266959
rect 148465 266931 148499 266959
rect 148527 266931 148561 266959
rect 148589 266931 148623 266959
rect 148651 266931 157437 266959
rect 157465 266931 157499 266959
rect 157527 266931 157561 266959
rect 157589 266931 157623 266959
rect 157651 266931 166437 266959
rect 166465 266931 166499 266959
rect 166527 266931 166561 266959
rect 166589 266931 166623 266959
rect 166651 266931 175437 266959
rect 175465 266931 175499 266959
rect 175527 266931 175561 266959
rect 175589 266931 175623 266959
rect 175651 266931 184437 266959
rect 184465 266931 184499 266959
rect 184527 266931 184561 266959
rect 184589 266931 184623 266959
rect 184651 266931 193437 266959
rect 193465 266931 193499 266959
rect 193527 266931 193561 266959
rect 193589 266931 193623 266959
rect 193651 266931 202437 266959
rect 202465 266931 202499 266959
rect 202527 266931 202561 266959
rect 202589 266931 202623 266959
rect 202651 266931 211437 266959
rect 211465 266931 211499 266959
rect 211527 266931 211561 266959
rect 211589 266931 211623 266959
rect 211651 266931 220437 266959
rect 220465 266931 220499 266959
rect 220527 266931 220561 266959
rect 220589 266931 220623 266959
rect 220651 266931 229437 266959
rect 229465 266931 229499 266959
rect 229527 266931 229561 266959
rect 229589 266931 229623 266959
rect 229651 266931 238437 266959
rect 238465 266931 238499 266959
rect 238527 266931 238561 266959
rect 238589 266931 238623 266959
rect 238651 266931 247437 266959
rect 247465 266931 247499 266959
rect 247527 266931 247561 266959
rect 247589 266931 247623 266959
rect 247651 266931 256437 266959
rect 256465 266931 256499 266959
rect 256527 266931 256561 266959
rect 256589 266931 256623 266959
rect 256651 266931 265437 266959
rect 265465 266931 265499 266959
rect 265527 266931 265561 266959
rect 265589 266931 265623 266959
rect 265651 266931 274437 266959
rect 274465 266931 274499 266959
rect 274527 266931 274561 266959
rect 274589 266931 274623 266959
rect 274651 266931 283437 266959
rect 283465 266931 283499 266959
rect 283527 266931 283561 266959
rect 283589 266931 283623 266959
rect 283651 266931 292437 266959
rect 292465 266931 292499 266959
rect 292527 266931 292561 266959
rect 292589 266931 292623 266959
rect 292651 266931 299736 266959
rect 299764 266931 299798 266959
rect 299826 266931 299860 266959
rect 299888 266931 299922 266959
rect 299950 266931 299998 266959
rect -6 266897 299998 266931
rect -6 266869 42 266897
rect 70 266869 104 266897
rect 132 266869 166 266897
rect 194 266869 228 266897
rect 256 266869 4437 266897
rect 4465 266869 4499 266897
rect 4527 266869 4561 266897
rect 4589 266869 4623 266897
rect 4651 266869 13437 266897
rect 13465 266869 13499 266897
rect 13527 266869 13561 266897
rect 13589 266869 13623 266897
rect 13651 266869 22437 266897
rect 22465 266869 22499 266897
rect 22527 266869 22561 266897
rect 22589 266869 22623 266897
rect 22651 266869 31437 266897
rect 31465 266869 31499 266897
rect 31527 266869 31561 266897
rect 31589 266869 31623 266897
rect 31651 266869 40437 266897
rect 40465 266869 40499 266897
rect 40527 266869 40561 266897
rect 40589 266869 40623 266897
rect 40651 266869 49437 266897
rect 49465 266869 49499 266897
rect 49527 266869 49561 266897
rect 49589 266869 49623 266897
rect 49651 266869 58437 266897
rect 58465 266869 58499 266897
rect 58527 266869 58561 266897
rect 58589 266869 58623 266897
rect 58651 266869 67437 266897
rect 67465 266869 67499 266897
rect 67527 266869 67561 266897
rect 67589 266869 67623 266897
rect 67651 266869 76437 266897
rect 76465 266869 76499 266897
rect 76527 266869 76561 266897
rect 76589 266869 76623 266897
rect 76651 266869 85437 266897
rect 85465 266869 85499 266897
rect 85527 266869 85561 266897
rect 85589 266869 85623 266897
rect 85651 266869 94437 266897
rect 94465 266869 94499 266897
rect 94527 266869 94561 266897
rect 94589 266869 94623 266897
rect 94651 266869 103437 266897
rect 103465 266869 103499 266897
rect 103527 266869 103561 266897
rect 103589 266869 103623 266897
rect 103651 266869 112437 266897
rect 112465 266869 112499 266897
rect 112527 266869 112561 266897
rect 112589 266869 112623 266897
rect 112651 266869 121437 266897
rect 121465 266869 121499 266897
rect 121527 266869 121561 266897
rect 121589 266869 121623 266897
rect 121651 266869 130437 266897
rect 130465 266869 130499 266897
rect 130527 266869 130561 266897
rect 130589 266869 130623 266897
rect 130651 266869 139437 266897
rect 139465 266869 139499 266897
rect 139527 266869 139561 266897
rect 139589 266869 139623 266897
rect 139651 266869 148437 266897
rect 148465 266869 148499 266897
rect 148527 266869 148561 266897
rect 148589 266869 148623 266897
rect 148651 266869 157437 266897
rect 157465 266869 157499 266897
rect 157527 266869 157561 266897
rect 157589 266869 157623 266897
rect 157651 266869 166437 266897
rect 166465 266869 166499 266897
rect 166527 266869 166561 266897
rect 166589 266869 166623 266897
rect 166651 266869 175437 266897
rect 175465 266869 175499 266897
rect 175527 266869 175561 266897
rect 175589 266869 175623 266897
rect 175651 266869 184437 266897
rect 184465 266869 184499 266897
rect 184527 266869 184561 266897
rect 184589 266869 184623 266897
rect 184651 266869 193437 266897
rect 193465 266869 193499 266897
rect 193527 266869 193561 266897
rect 193589 266869 193623 266897
rect 193651 266869 202437 266897
rect 202465 266869 202499 266897
rect 202527 266869 202561 266897
rect 202589 266869 202623 266897
rect 202651 266869 211437 266897
rect 211465 266869 211499 266897
rect 211527 266869 211561 266897
rect 211589 266869 211623 266897
rect 211651 266869 220437 266897
rect 220465 266869 220499 266897
rect 220527 266869 220561 266897
rect 220589 266869 220623 266897
rect 220651 266869 229437 266897
rect 229465 266869 229499 266897
rect 229527 266869 229561 266897
rect 229589 266869 229623 266897
rect 229651 266869 238437 266897
rect 238465 266869 238499 266897
rect 238527 266869 238561 266897
rect 238589 266869 238623 266897
rect 238651 266869 247437 266897
rect 247465 266869 247499 266897
rect 247527 266869 247561 266897
rect 247589 266869 247623 266897
rect 247651 266869 256437 266897
rect 256465 266869 256499 266897
rect 256527 266869 256561 266897
rect 256589 266869 256623 266897
rect 256651 266869 265437 266897
rect 265465 266869 265499 266897
rect 265527 266869 265561 266897
rect 265589 266869 265623 266897
rect 265651 266869 274437 266897
rect 274465 266869 274499 266897
rect 274527 266869 274561 266897
rect 274589 266869 274623 266897
rect 274651 266869 283437 266897
rect 283465 266869 283499 266897
rect 283527 266869 283561 266897
rect 283589 266869 283623 266897
rect 283651 266869 292437 266897
rect 292465 266869 292499 266897
rect 292527 266869 292561 266897
rect 292589 266869 292623 266897
rect 292651 266869 299736 266897
rect 299764 266869 299798 266897
rect 299826 266869 299860 266897
rect 299888 266869 299922 266897
rect 299950 266869 299998 266897
rect -6 266835 299998 266869
rect -6 266807 42 266835
rect 70 266807 104 266835
rect 132 266807 166 266835
rect 194 266807 228 266835
rect 256 266807 4437 266835
rect 4465 266807 4499 266835
rect 4527 266807 4561 266835
rect 4589 266807 4623 266835
rect 4651 266807 13437 266835
rect 13465 266807 13499 266835
rect 13527 266807 13561 266835
rect 13589 266807 13623 266835
rect 13651 266807 22437 266835
rect 22465 266807 22499 266835
rect 22527 266807 22561 266835
rect 22589 266807 22623 266835
rect 22651 266807 31437 266835
rect 31465 266807 31499 266835
rect 31527 266807 31561 266835
rect 31589 266807 31623 266835
rect 31651 266807 40437 266835
rect 40465 266807 40499 266835
rect 40527 266807 40561 266835
rect 40589 266807 40623 266835
rect 40651 266807 49437 266835
rect 49465 266807 49499 266835
rect 49527 266807 49561 266835
rect 49589 266807 49623 266835
rect 49651 266807 58437 266835
rect 58465 266807 58499 266835
rect 58527 266807 58561 266835
rect 58589 266807 58623 266835
rect 58651 266807 67437 266835
rect 67465 266807 67499 266835
rect 67527 266807 67561 266835
rect 67589 266807 67623 266835
rect 67651 266807 76437 266835
rect 76465 266807 76499 266835
rect 76527 266807 76561 266835
rect 76589 266807 76623 266835
rect 76651 266807 85437 266835
rect 85465 266807 85499 266835
rect 85527 266807 85561 266835
rect 85589 266807 85623 266835
rect 85651 266807 94437 266835
rect 94465 266807 94499 266835
rect 94527 266807 94561 266835
rect 94589 266807 94623 266835
rect 94651 266807 103437 266835
rect 103465 266807 103499 266835
rect 103527 266807 103561 266835
rect 103589 266807 103623 266835
rect 103651 266807 112437 266835
rect 112465 266807 112499 266835
rect 112527 266807 112561 266835
rect 112589 266807 112623 266835
rect 112651 266807 121437 266835
rect 121465 266807 121499 266835
rect 121527 266807 121561 266835
rect 121589 266807 121623 266835
rect 121651 266807 130437 266835
rect 130465 266807 130499 266835
rect 130527 266807 130561 266835
rect 130589 266807 130623 266835
rect 130651 266807 139437 266835
rect 139465 266807 139499 266835
rect 139527 266807 139561 266835
rect 139589 266807 139623 266835
rect 139651 266807 148437 266835
rect 148465 266807 148499 266835
rect 148527 266807 148561 266835
rect 148589 266807 148623 266835
rect 148651 266807 157437 266835
rect 157465 266807 157499 266835
rect 157527 266807 157561 266835
rect 157589 266807 157623 266835
rect 157651 266807 166437 266835
rect 166465 266807 166499 266835
rect 166527 266807 166561 266835
rect 166589 266807 166623 266835
rect 166651 266807 175437 266835
rect 175465 266807 175499 266835
rect 175527 266807 175561 266835
rect 175589 266807 175623 266835
rect 175651 266807 184437 266835
rect 184465 266807 184499 266835
rect 184527 266807 184561 266835
rect 184589 266807 184623 266835
rect 184651 266807 193437 266835
rect 193465 266807 193499 266835
rect 193527 266807 193561 266835
rect 193589 266807 193623 266835
rect 193651 266807 202437 266835
rect 202465 266807 202499 266835
rect 202527 266807 202561 266835
rect 202589 266807 202623 266835
rect 202651 266807 211437 266835
rect 211465 266807 211499 266835
rect 211527 266807 211561 266835
rect 211589 266807 211623 266835
rect 211651 266807 220437 266835
rect 220465 266807 220499 266835
rect 220527 266807 220561 266835
rect 220589 266807 220623 266835
rect 220651 266807 229437 266835
rect 229465 266807 229499 266835
rect 229527 266807 229561 266835
rect 229589 266807 229623 266835
rect 229651 266807 238437 266835
rect 238465 266807 238499 266835
rect 238527 266807 238561 266835
rect 238589 266807 238623 266835
rect 238651 266807 247437 266835
rect 247465 266807 247499 266835
rect 247527 266807 247561 266835
rect 247589 266807 247623 266835
rect 247651 266807 256437 266835
rect 256465 266807 256499 266835
rect 256527 266807 256561 266835
rect 256589 266807 256623 266835
rect 256651 266807 265437 266835
rect 265465 266807 265499 266835
rect 265527 266807 265561 266835
rect 265589 266807 265623 266835
rect 265651 266807 274437 266835
rect 274465 266807 274499 266835
rect 274527 266807 274561 266835
rect 274589 266807 274623 266835
rect 274651 266807 283437 266835
rect 283465 266807 283499 266835
rect 283527 266807 283561 266835
rect 283589 266807 283623 266835
rect 283651 266807 292437 266835
rect 292465 266807 292499 266835
rect 292527 266807 292561 266835
rect 292589 266807 292623 266835
rect 292651 266807 299736 266835
rect 299764 266807 299798 266835
rect 299826 266807 299860 266835
rect 299888 266807 299922 266835
rect 299950 266807 299998 266835
rect -6 266773 299998 266807
rect -6 266745 42 266773
rect 70 266745 104 266773
rect 132 266745 166 266773
rect 194 266745 228 266773
rect 256 266745 4437 266773
rect 4465 266745 4499 266773
rect 4527 266745 4561 266773
rect 4589 266745 4623 266773
rect 4651 266745 13437 266773
rect 13465 266745 13499 266773
rect 13527 266745 13561 266773
rect 13589 266745 13623 266773
rect 13651 266745 22437 266773
rect 22465 266745 22499 266773
rect 22527 266745 22561 266773
rect 22589 266745 22623 266773
rect 22651 266745 31437 266773
rect 31465 266745 31499 266773
rect 31527 266745 31561 266773
rect 31589 266745 31623 266773
rect 31651 266745 40437 266773
rect 40465 266745 40499 266773
rect 40527 266745 40561 266773
rect 40589 266745 40623 266773
rect 40651 266745 49437 266773
rect 49465 266745 49499 266773
rect 49527 266745 49561 266773
rect 49589 266745 49623 266773
rect 49651 266745 58437 266773
rect 58465 266745 58499 266773
rect 58527 266745 58561 266773
rect 58589 266745 58623 266773
rect 58651 266745 67437 266773
rect 67465 266745 67499 266773
rect 67527 266745 67561 266773
rect 67589 266745 67623 266773
rect 67651 266745 76437 266773
rect 76465 266745 76499 266773
rect 76527 266745 76561 266773
rect 76589 266745 76623 266773
rect 76651 266745 85437 266773
rect 85465 266745 85499 266773
rect 85527 266745 85561 266773
rect 85589 266745 85623 266773
rect 85651 266745 94437 266773
rect 94465 266745 94499 266773
rect 94527 266745 94561 266773
rect 94589 266745 94623 266773
rect 94651 266745 103437 266773
rect 103465 266745 103499 266773
rect 103527 266745 103561 266773
rect 103589 266745 103623 266773
rect 103651 266745 112437 266773
rect 112465 266745 112499 266773
rect 112527 266745 112561 266773
rect 112589 266745 112623 266773
rect 112651 266745 121437 266773
rect 121465 266745 121499 266773
rect 121527 266745 121561 266773
rect 121589 266745 121623 266773
rect 121651 266745 130437 266773
rect 130465 266745 130499 266773
rect 130527 266745 130561 266773
rect 130589 266745 130623 266773
rect 130651 266745 139437 266773
rect 139465 266745 139499 266773
rect 139527 266745 139561 266773
rect 139589 266745 139623 266773
rect 139651 266745 148437 266773
rect 148465 266745 148499 266773
rect 148527 266745 148561 266773
rect 148589 266745 148623 266773
rect 148651 266745 157437 266773
rect 157465 266745 157499 266773
rect 157527 266745 157561 266773
rect 157589 266745 157623 266773
rect 157651 266745 166437 266773
rect 166465 266745 166499 266773
rect 166527 266745 166561 266773
rect 166589 266745 166623 266773
rect 166651 266745 175437 266773
rect 175465 266745 175499 266773
rect 175527 266745 175561 266773
rect 175589 266745 175623 266773
rect 175651 266745 184437 266773
rect 184465 266745 184499 266773
rect 184527 266745 184561 266773
rect 184589 266745 184623 266773
rect 184651 266745 193437 266773
rect 193465 266745 193499 266773
rect 193527 266745 193561 266773
rect 193589 266745 193623 266773
rect 193651 266745 202437 266773
rect 202465 266745 202499 266773
rect 202527 266745 202561 266773
rect 202589 266745 202623 266773
rect 202651 266745 211437 266773
rect 211465 266745 211499 266773
rect 211527 266745 211561 266773
rect 211589 266745 211623 266773
rect 211651 266745 220437 266773
rect 220465 266745 220499 266773
rect 220527 266745 220561 266773
rect 220589 266745 220623 266773
rect 220651 266745 229437 266773
rect 229465 266745 229499 266773
rect 229527 266745 229561 266773
rect 229589 266745 229623 266773
rect 229651 266745 238437 266773
rect 238465 266745 238499 266773
rect 238527 266745 238561 266773
rect 238589 266745 238623 266773
rect 238651 266745 247437 266773
rect 247465 266745 247499 266773
rect 247527 266745 247561 266773
rect 247589 266745 247623 266773
rect 247651 266745 256437 266773
rect 256465 266745 256499 266773
rect 256527 266745 256561 266773
rect 256589 266745 256623 266773
rect 256651 266745 265437 266773
rect 265465 266745 265499 266773
rect 265527 266745 265561 266773
rect 265589 266745 265623 266773
rect 265651 266745 274437 266773
rect 274465 266745 274499 266773
rect 274527 266745 274561 266773
rect 274589 266745 274623 266773
rect 274651 266745 283437 266773
rect 283465 266745 283499 266773
rect 283527 266745 283561 266773
rect 283589 266745 283623 266773
rect 283651 266745 292437 266773
rect 292465 266745 292499 266773
rect 292527 266745 292561 266773
rect 292589 266745 292623 266773
rect 292651 266745 299736 266773
rect 299764 266745 299798 266773
rect 299826 266745 299860 266773
rect 299888 266745 299922 266773
rect 299950 266745 299998 266773
rect -6 266697 299998 266745
rect -6 263959 299998 264007
rect -6 263931 522 263959
rect 550 263931 584 263959
rect 612 263931 646 263959
rect 674 263931 708 263959
rect 736 263931 2577 263959
rect 2605 263931 2639 263959
rect 2667 263931 2701 263959
rect 2729 263931 2763 263959
rect 2791 263931 11577 263959
rect 11605 263931 11639 263959
rect 11667 263931 11701 263959
rect 11729 263931 11763 263959
rect 11791 263931 20577 263959
rect 20605 263931 20639 263959
rect 20667 263931 20701 263959
rect 20729 263931 20763 263959
rect 20791 263931 29577 263959
rect 29605 263931 29639 263959
rect 29667 263931 29701 263959
rect 29729 263931 29763 263959
rect 29791 263931 38577 263959
rect 38605 263931 38639 263959
rect 38667 263931 38701 263959
rect 38729 263931 38763 263959
rect 38791 263931 47577 263959
rect 47605 263931 47639 263959
rect 47667 263931 47701 263959
rect 47729 263931 47763 263959
rect 47791 263931 56577 263959
rect 56605 263931 56639 263959
rect 56667 263931 56701 263959
rect 56729 263931 56763 263959
rect 56791 263931 65577 263959
rect 65605 263931 65639 263959
rect 65667 263931 65701 263959
rect 65729 263931 65763 263959
rect 65791 263931 74577 263959
rect 74605 263931 74639 263959
rect 74667 263931 74701 263959
rect 74729 263931 74763 263959
rect 74791 263931 83577 263959
rect 83605 263931 83639 263959
rect 83667 263931 83701 263959
rect 83729 263931 83763 263959
rect 83791 263931 92577 263959
rect 92605 263931 92639 263959
rect 92667 263931 92701 263959
rect 92729 263931 92763 263959
rect 92791 263931 101577 263959
rect 101605 263931 101639 263959
rect 101667 263931 101701 263959
rect 101729 263931 101763 263959
rect 101791 263931 110577 263959
rect 110605 263931 110639 263959
rect 110667 263931 110701 263959
rect 110729 263931 110763 263959
rect 110791 263931 119577 263959
rect 119605 263931 119639 263959
rect 119667 263931 119701 263959
rect 119729 263931 119763 263959
rect 119791 263931 128577 263959
rect 128605 263931 128639 263959
rect 128667 263931 128701 263959
rect 128729 263931 128763 263959
rect 128791 263931 137577 263959
rect 137605 263931 137639 263959
rect 137667 263931 137701 263959
rect 137729 263931 137763 263959
rect 137791 263931 146577 263959
rect 146605 263931 146639 263959
rect 146667 263931 146701 263959
rect 146729 263931 146763 263959
rect 146791 263931 155577 263959
rect 155605 263931 155639 263959
rect 155667 263931 155701 263959
rect 155729 263931 155763 263959
rect 155791 263931 164577 263959
rect 164605 263931 164639 263959
rect 164667 263931 164701 263959
rect 164729 263931 164763 263959
rect 164791 263931 173577 263959
rect 173605 263931 173639 263959
rect 173667 263931 173701 263959
rect 173729 263931 173763 263959
rect 173791 263931 182577 263959
rect 182605 263931 182639 263959
rect 182667 263931 182701 263959
rect 182729 263931 182763 263959
rect 182791 263931 191577 263959
rect 191605 263931 191639 263959
rect 191667 263931 191701 263959
rect 191729 263931 191763 263959
rect 191791 263931 200577 263959
rect 200605 263931 200639 263959
rect 200667 263931 200701 263959
rect 200729 263931 200763 263959
rect 200791 263931 209577 263959
rect 209605 263931 209639 263959
rect 209667 263931 209701 263959
rect 209729 263931 209763 263959
rect 209791 263931 218577 263959
rect 218605 263931 218639 263959
rect 218667 263931 218701 263959
rect 218729 263931 218763 263959
rect 218791 263931 227577 263959
rect 227605 263931 227639 263959
rect 227667 263931 227701 263959
rect 227729 263931 227763 263959
rect 227791 263931 236577 263959
rect 236605 263931 236639 263959
rect 236667 263931 236701 263959
rect 236729 263931 236763 263959
rect 236791 263931 245577 263959
rect 245605 263931 245639 263959
rect 245667 263931 245701 263959
rect 245729 263931 245763 263959
rect 245791 263931 254577 263959
rect 254605 263931 254639 263959
rect 254667 263931 254701 263959
rect 254729 263931 254763 263959
rect 254791 263931 263577 263959
rect 263605 263931 263639 263959
rect 263667 263931 263701 263959
rect 263729 263931 263763 263959
rect 263791 263931 272577 263959
rect 272605 263931 272639 263959
rect 272667 263931 272701 263959
rect 272729 263931 272763 263959
rect 272791 263931 281577 263959
rect 281605 263931 281639 263959
rect 281667 263931 281701 263959
rect 281729 263931 281763 263959
rect 281791 263931 290577 263959
rect 290605 263931 290639 263959
rect 290667 263931 290701 263959
rect 290729 263931 290763 263959
rect 290791 263931 299256 263959
rect 299284 263931 299318 263959
rect 299346 263931 299380 263959
rect 299408 263931 299442 263959
rect 299470 263931 299998 263959
rect -6 263897 299998 263931
rect -6 263869 522 263897
rect 550 263869 584 263897
rect 612 263869 646 263897
rect 674 263869 708 263897
rect 736 263869 2577 263897
rect 2605 263869 2639 263897
rect 2667 263869 2701 263897
rect 2729 263869 2763 263897
rect 2791 263869 11577 263897
rect 11605 263869 11639 263897
rect 11667 263869 11701 263897
rect 11729 263869 11763 263897
rect 11791 263869 20577 263897
rect 20605 263869 20639 263897
rect 20667 263869 20701 263897
rect 20729 263869 20763 263897
rect 20791 263869 29577 263897
rect 29605 263869 29639 263897
rect 29667 263869 29701 263897
rect 29729 263869 29763 263897
rect 29791 263869 38577 263897
rect 38605 263869 38639 263897
rect 38667 263869 38701 263897
rect 38729 263869 38763 263897
rect 38791 263869 47577 263897
rect 47605 263869 47639 263897
rect 47667 263869 47701 263897
rect 47729 263869 47763 263897
rect 47791 263869 56577 263897
rect 56605 263869 56639 263897
rect 56667 263869 56701 263897
rect 56729 263869 56763 263897
rect 56791 263869 65577 263897
rect 65605 263869 65639 263897
rect 65667 263869 65701 263897
rect 65729 263869 65763 263897
rect 65791 263869 74577 263897
rect 74605 263869 74639 263897
rect 74667 263869 74701 263897
rect 74729 263869 74763 263897
rect 74791 263869 83577 263897
rect 83605 263869 83639 263897
rect 83667 263869 83701 263897
rect 83729 263869 83763 263897
rect 83791 263869 92577 263897
rect 92605 263869 92639 263897
rect 92667 263869 92701 263897
rect 92729 263869 92763 263897
rect 92791 263869 101577 263897
rect 101605 263869 101639 263897
rect 101667 263869 101701 263897
rect 101729 263869 101763 263897
rect 101791 263869 110577 263897
rect 110605 263869 110639 263897
rect 110667 263869 110701 263897
rect 110729 263869 110763 263897
rect 110791 263869 119577 263897
rect 119605 263869 119639 263897
rect 119667 263869 119701 263897
rect 119729 263869 119763 263897
rect 119791 263869 128577 263897
rect 128605 263869 128639 263897
rect 128667 263869 128701 263897
rect 128729 263869 128763 263897
rect 128791 263869 137577 263897
rect 137605 263869 137639 263897
rect 137667 263869 137701 263897
rect 137729 263869 137763 263897
rect 137791 263869 146577 263897
rect 146605 263869 146639 263897
rect 146667 263869 146701 263897
rect 146729 263869 146763 263897
rect 146791 263869 155577 263897
rect 155605 263869 155639 263897
rect 155667 263869 155701 263897
rect 155729 263869 155763 263897
rect 155791 263869 164577 263897
rect 164605 263869 164639 263897
rect 164667 263869 164701 263897
rect 164729 263869 164763 263897
rect 164791 263869 173577 263897
rect 173605 263869 173639 263897
rect 173667 263869 173701 263897
rect 173729 263869 173763 263897
rect 173791 263869 182577 263897
rect 182605 263869 182639 263897
rect 182667 263869 182701 263897
rect 182729 263869 182763 263897
rect 182791 263869 191577 263897
rect 191605 263869 191639 263897
rect 191667 263869 191701 263897
rect 191729 263869 191763 263897
rect 191791 263869 200577 263897
rect 200605 263869 200639 263897
rect 200667 263869 200701 263897
rect 200729 263869 200763 263897
rect 200791 263869 209577 263897
rect 209605 263869 209639 263897
rect 209667 263869 209701 263897
rect 209729 263869 209763 263897
rect 209791 263869 218577 263897
rect 218605 263869 218639 263897
rect 218667 263869 218701 263897
rect 218729 263869 218763 263897
rect 218791 263869 227577 263897
rect 227605 263869 227639 263897
rect 227667 263869 227701 263897
rect 227729 263869 227763 263897
rect 227791 263869 236577 263897
rect 236605 263869 236639 263897
rect 236667 263869 236701 263897
rect 236729 263869 236763 263897
rect 236791 263869 245577 263897
rect 245605 263869 245639 263897
rect 245667 263869 245701 263897
rect 245729 263869 245763 263897
rect 245791 263869 254577 263897
rect 254605 263869 254639 263897
rect 254667 263869 254701 263897
rect 254729 263869 254763 263897
rect 254791 263869 263577 263897
rect 263605 263869 263639 263897
rect 263667 263869 263701 263897
rect 263729 263869 263763 263897
rect 263791 263869 272577 263897
rect 272605 263869 272639 263897
rect 272667 263869 272701 263897
rect 272729 263869 272763 263897
rect 272791 263869 281577 263897
rect 281605 263869 281639 263897
rect 281667 263869 281701 263897
rect 281729 263869 281763 263897
rect 281791 263869 290577 263897
rect 290605 263869 290639 263897
rect 290667 263869 290701 263897
rect 290729 263869 290763 263897
rect 290791 263869 299256 263897
rect 299284 263869 299318 263897
rect 299346 263869 299380 263897
rect 299408 263869 299442 263897
rect 299470 263869 299998 263897
rect -6 263835 299998 263869
rect -6 263807 522 263835
rect 550 263807 584 263835
rect 612 263807 646 263835
rect 674 263807 708 263835
rect 736 263807 2577 263835
rect 2605 263807 2639 263835
rect 2667 263807 2701 263835
rect 2729 263807 2763 263835
rect 2791 263807 11577 263835
rect 11605 263807 11639 263835
rect 11667 263807 11701 263835
rect 11729 263807 11763 263835
rect 11791 263807 20577 263835
rect 20605 263807 20639 263835
rect 20667 263807 20701 263835
rect 20729 263807 20763 263835
rect 20791 263807 29577 263835
rect 29605 263807 29639 263835
rect 29667 263807 29701 263835
rect 29729 263807 29763 263835
rect 29791 263807 38577 263835
rect 38605 263807 38639 263835
rect 38667 263807 38701 263835
rect 38729 263807 38763 263835
rect 38791 263807 47577 263835
rect 47605 263807 47639 263835
rect 47667 263807 47701 263835
rect 47729 263807 47763 263835
rect 47791 263807 56577 263835
rect 56605 263807 56639 263835
rect 56667 263807 56701 263835
rect 56729 263807 56763 263835
rect 56791 263807 65577 263835
rect 65605 263807 65639 263835
rect 65667 263807 65701 263835
rect 65729 263807 65763 263835
rect 65791 263807 74577 263835
rect 74605 263807 74639 263835
rect 74667 263807 74701 263835
rect 74729 263807 74763 263835
rect 74791 263807 83577 263835
rect 83605 263807 83639 263835
rect 83667 263807 83701 263835
rect 83729 263807 83763 263835
rect 83791 263807 92577 263835
rect 92605 263807 92639 263835
rect 92667 263807 92701 263835
rect 92729 263807 92763 263835
rect 92791 263807 101577 263835
rect 101605 263807 101639 263835
rect 101667 263807 101701 263835
rect 101729 263807 101763 263835
rect 101791 263807 110577 263835
rect 110605 263807 110639 263835
rect 110667 263807 110701 263835
rect 110729 263807 110763 263835
rect 110791 263807 119577 263835
rect 119605 263807 119639 263835
rect 119667 263807 119701 263835
rect 119729 263807 119763 263835
rect 119791 263807 128577 263835
rect 128605 263807 128639 263835
rect 128667 263807 128701 263835
rect 128729 263807 128763 263835
rect 128791 263807 137577 263835
rect 137605 263807 137639 263835
rect 137667 263807 137701 263835
rect 137729 263807 137763 263835
rect 137791 263807 146577 263835
rect 146605 263807 146639 263835
rect 146667 263807 146701 263835
rect 146729 263807 146763 263835
rect 146791 263807 155577 263835
rect 155605 263807 155639 263835
rect 155667 263807 155701 263835
rect 155729 263807 155763 263835
rect 155791 263807 164577 263835
rect 164605 263807 164639 263835
rect 164667 263807 164701 263835
rect 164729 263807 164763 263835
rect 164791 263807 173577 263835
rect 173605 263807 173639 263835
rect 173667 263807 173701 263835
rect 173729 263807 173763 263835
rect 173791 263807 182577 263835
rect 182605 263807 182639 263835
rect 182667 263807 182701 263835
rect 182729 263807 182763 263835
rect 182791 263807 191577 263835
rect 191605 263807 191639 263835
rect 191667 263807 191701 263835
rect 191729 263807 191763 263835
rect 191791 263807 200577 263835
rect 200605 263807 200639 263835
rect 200667 263807 200701 263835
rect 200729 263807 200763 263835
rect 200791 263807 209577 263835
rect 209605 263807 209639 263835
rect 209667 263807 209701 263835
rect 209729 263807 209763 263835
rect 209791 263807 218577 263835
rect 218605 263807 218639 263835
rect 218667 263807 218701 263835
rect 218729 263807 218763 263835
rect 218791 263807 227577 263835
rect 227605 263807 227639 263835
rect 227667 263807 227701 263835
rect 227729 263807 227763 263835
rect 227791 263807 236577 263835
rect 236605 263807 236639 263835
rect 236667 263807 236701 263835
rect 236729 263807 236763 263835
rect 236791 263807 245577 263835
rect 245605 263807 245639 263835
rect 245667 263807 245701 263835
rect 245729 263807 245763 263835
rect 245791 263807 254577 263835
rect 254605 263807 254639 263835
rect 254667 263807 254701 263835
rect 254729 263807 254763 263835
rect 254791 263807 263577 263835
rect 263605 263807 263639 263835
rect 263667 263807 263701 263835
rect 263729 263807 263763 263835
rect 263791 263807 272577 263835
rect 272605 263807 272639 263835
rect 272667 263807 272701 263835
rect 272729 263807 272763 263835
rect 272791 263807 281577 263835
rect 281605 263807 281639 263835
rect 281667 263807 281701 263835
rect 281729 263807 281763 263835
rect 281791 263807 290577 263835
rect 290605 263807 290639 263835
rect 290667 263807 290701 263835
rect 290729 263807 290763 263835
rect 290791 263807 299256 263835
rect 299284 263807 299318 263835
rect 299346 263807 299380 263835
rect 299408 263807 299442 263835
rect 299470 263807 299998 263835
rect -6 263773 299998 263807
rect -6 263745 522 263773
rect 550 263745 584 263773
rect 612 263745 646 263773
rect 674 263745 708 263773
rect 736 263745 2577 263773
rect 2605 263745 2639 263773
rect 2667 263745 2701 263773
rect 2729 263745 2763 263773
rect 2791 263745 11577 263773
rect 11605 263745 11639 263773
rect 11667 263745 11701 263773
rect 11729 263745 11763 263773
rect 11791 263745 20577 263773
rect 20605 263745 20639 263773
rect 20667 263745 20701 263773
rect 20729 263745 20763 263773
rect 20791 263745 29577 263773
rect 29605 263745 29639 263773
rect 29667 263745 29701 263773
rect 29729 263745 29763 263773
rect 29791 263745 38577 263773
rect 38605 263745 38639 263773
rect 38667 263745 38701 263773
rect 38729 263745 38763 263773
rect 38791 263745 47577 263773
rect 47605 263745 47639 263773
rect 47667 263745 47701 263773
rect 47729 263745 47763 263773
rect 47791 263745 56577 263773
rect 56605 263745 56639 263773
rect 56667 263745 56701 263773
rect 56729 263745 56763 263773
rect 56791 263745 65577 263773
rect 65605 263745 65639 263773
rect 65667 263745 65701 263773
rect 65729 263745 65763 263773
rect 65791 263745 74577 263773
rect 74605 263745 74639 263773
rect 74667 263745 74701 263773
rect 74729 263745 74763 263773
rect 74791 263745 83577 263773
rect 83605 263745 83639 263773
rect 83667 263745 83701 263773
rect 83729 263745 83763 263773
rect 83791 263745 92577 263773
rect 92605 263745 92639 263773
rect 92667 263745 92701 263773
rect 92729 263745 92763 263773
rect 92791 263745 101577 263773
rect 101605 263745 101639 263773
rect 101667 263745 101701 263773
rect 101729 263745 101763 263773
rect 101791 263745 110577 263773
rect 110605 263745 110639 263773
rect 110667 263745 110701 263773
rect 110729 263745 110763 263773
rect 110791 263745 119577 263773
rect 119605 263745 119639 263773
rect 119667 263745 119701 263773
rect 119729 263745 119763 263773
rect 119791 263745 128577 263773
rect 128605 263745 128639 263773
rect 128667 263745 128701 263773
rect 128729 263745 128763 263773
rect 128791 263745 137577 263773
rect 137605 263745 137639 263773
rect 137667 263745 137701 263773
rect 137729 263745 137763 263773
rect 137791 263745 146577 263773
rect 146605 263745 146639 263773
rect 146667 263745 146701 263773
rect 146729 263745 146763 263773
rect 146791 263745 155577 263773
rect 155605 263745 155639 263773
rect 155667 263745 155701 263773
rect 155729 263745 155763 263773
rect 155791 263745 164577 263773
rect 164605 263745 164639 263773
rect 164667 263745 164701 263773
rect 164729 263745 164763 263773
rect 164791 263745 173577 263773
rect 173605 263745 173639 263773
rect 173667 263745 173701 263773
rect 173729 263745 173763 263773
rect 173791 263745 182577 263773
rect 182605 263745 182639 263773
rect 182667 263745 182701 263773
rect 182729 263745 182763 263773
rect 182791 263745 191577 263773
rect 191605 263745 191639 263773
rect 191667 263745 191701 263773
rect 191729 263745 191763 263773
rect 191791 263745 200577 263773
rect 200605 263745 200639 263773
rect 200667 263745 200701 263773
rect 200729 263745 200763 263773
rect 200791 263745 209577 263773
rect 209605 263745 209639 263773
rect 209667 263745 209701 263773
rect 209729 263745 209763 263773
rect 209791 263745 218577 263773
rect 218605 263745 218639 263773
rect 218667 263745 218701 263773
rect 218729 263745 218763 263773
rect 218791 263745 227577 263773
rect 227605 263745 227639 263773
rect 227667 263745 227701 263773
rect 227729 263745 227763 263773
rect 227791 263745 236577 263773
rect 236605 263745 236639 263773
rect 236667 263745 236701 263773
rect 236729 263745 236763 263773
rect 236791 263745 245577 263773
rect 245605 263745 245639 263773
rect 245667 263745 245701 263773
rect 245729 263745 245763 263773
rect 245791 263745 254577 263773
rect 254605 263745 254639 263773
rect 254667 263745 254701 263773
rect 254729 263745 254763 263773
rect 254791 263745 263577 263773
rect 263605 263745 263639 263773
rect 263667 263745 263701 263773
rect 263729 263745 263763 263773
rect 263791 263745 272577 263773
rect 272605 263745 272639 263773
rect 272667 263745 272701 263773
rect 272729 263745 272763 263773
rect 272791 263745 281577 263773
rect 281605 263745 281639 263773
rect 281667 263745 281701 263773
rect 281729 263745 281763 263773
rect 281791 263745 290577 263773
rect 290605 263745 290639 263773
rect 290667 263745 290701 263773
rect 290729 263745 290763 263773
rect 290791 263745 299256 263773
rect 299284 263745 299318 263773
rect 299346 263745 299380 263773
rect 299408 263745 299442 263773
rect 299470 263745 299998 263773
rect -6 263697 299998 263745
rect -6 257959 299998 258007
rect -6 257931 42 257959
rect 70 257931 104 257959
rect 132 257931 166 257959
rect 194 257931 228 257959
rect 256 257931 4437 257959
rect 4465 257931 4499 257959
rect 4527 257931 4561 257959
rect 4589 257931 4623 257959
rect 4651 257931 13437 257959
rect 13465 257931 13499 257959
rect 13527 257931 13561 257959
rect 13589 257931 13623 257959
rect 13651 257931 22437 257959
rect 22465 257931 22499 257959
rect 22527 257931 22561 257959
rect 22589 257931 22623 257959
rect 22651 257931 31437 257959
rect 31465 257931 31499 257959
rect 31527 257931 31561 257959
rect 31589 257931 31623 257959
rect 31651 257931 40437 257959
rect 40465 257931 40499 257959
rect 40527 257931 40561 257959
rect 40589 257931 40623 257959
rect 40651 257931 49437 257959
rect 49465 257931 49499 257959
rect 49527 257931 49561 257959
rect 49589 257931 49623 257959
rect 49651 257931 58437 257959
rect 58465 257931 58499 257959
rect 58527 257931 58561 257959
rect 58589 257931 58623 257959
rect 58651 257931 67437 257959
rect 67465 257931 67499 257959
rect 67527 257931 67561 257959
rect 67589 257931 67623 257959
rect 67651 257931 76437 257959
rect 76465 257931 76499 257959
rect 76527 257931 76561 257959
rect 76589 257931 76623 257959
rect 76651 257931 85437 257959
rect 85465 257931 85499 257959
rect 85527 257931 85561 257959
rect 85589 257931 85623 257959
rect 85651 257931 94437 257959
rect 94465 257931 94499 257959
rect 94527 257931 94561 257959
rect 94589 257931 94623 257959
rect 94651 257931 103437 257959
rect 103465 257931 103499 257959
rect 103527 257931 103561 257959
rect 103589 257931 103623 257959
rect 103651 257931 112437 257959
rect 112465 257931 112499 257959
rect 112527 257931 112561 257959
rect 112589 257931 112623 257959
rect 112651 257931 121437 257959
rect 121465 257931 121499 257959
rect 121527 257931 121561 257959
rect 121589 257931 121623 257959
rect 121651 257931 130437 257959
rect 130465 257931 130499 257959
rect 130527 257931 130561 257959
rect 130589 257931 130623 257959
rect 130651 257931 139437 257959
rect 139465 257931 139499 257959
rect 139527 257931 139561 257959
rect 139589 257931 139623 257959
rect 139651 257931 148437 257959
rect 148465 257931 148499 257959
rect 148527 257931 148561 257959
rect 148589 257931 148623 257959
rect 148651 257931 157437 257959
rect 157465 257931 157499 257959
rect 157527 257931 157561 257959
rect 157589 257931 157623 257959
rect 157651 257931 166437 257959
rect 166465 257931 166499 257959
rect 166527 257931 166561 257959
rect 166589 257931 166623 257959
rect 166651 257931 175437 257959
rect 175465 257931 175499 257959
rect 175527 257931 175561 257959
rect 175589 257931 175623 257959
rect 175651 257931 184437 257959
rect 184465 257931 184499 257959
rect 184527 257931 184561 257959
rect 184589 257931 184623 257959
rect 184651 257931 193437 257959
rect 193465 257931 193499 257959
rect 193527 257931 193561 257959
rect 193589 257931 193623 257959
rect 193651 257931 202437 257959
rect 202465 257931 202499 257959
rect 202527 257931 202561 257959
rect 202589 257931 202623 257959
rect 202651 257931 211437 257959
rect 211465 257931 211499 257959
rect 211527 257931 211561 257959
rect 211589 257931 211623 257959
rect 211651 257931 220437 257959
rect 220465 257931 220499 257959
rect 220527 257931 220561 257959
rect 220589 257931 220623 257959
rect 220651 257931 229437 257959
rect 229465 257931 229499 257959
rect 229527 257931 229561 257959
rect 229589 257931 229623 257959
rect 229651 257931 238437 257959
rect 238465 257931 238499 257959
rect 238527 257931 238561 257959
rect 238589 257931 238623 257959
rect 238651 257931 247437 257959
rect 247465 257931 247499 257959
rect 247527 257931 247561 257959
rect 247589 257931 247623 257959
rect 247651 257931 256437 257959
rect 256465 257931 256499 257959
rect 256527 257931 256561 257959
rect 256589 257931 256623 257959
rect 256651 257931 265437 257959
rect 265465 257931 265499 257959
rect 265527 257931 265561 257959
rect 265589 257931 265623 257959
rect 265651 257931 274437 257959
rect 274465 257931 274499 257959
rect 274527 257931 274561 257959
rect 274589 257931 274623 257959
rect 274651 257931 283437 257959
rect 283465 257931 283499 257959
rect 283527 257931 283561 257959
rect 283589 257931 283623 257959
rect 283651 257931 292437 257959
rect 292465 257931 292499 257959
rect 292527 257931 292561 257959
rect 292589 257931 292623 257959
rect 292651 257931 299736 257959
rect 299764 257931 299798 257959
rect 299826 257931 299860 257959
rect 299888 257931 299922 257959
rect 299950 257931 299998 257959
rect -6 257897 299998 257931
rect -6 257869 42 257897
rect 70 257869 104 257897
rect 132 257869 166 257897
rect 194 257869 228 257897
rect 256 257869 4437 257897
rect 4465 257869 4499 257897
rect 4527 257869 4561 257897
rect 4589 257869 4623 257897
rect 4651 257869 13437 257897
rect 13465 257869 13499 257897
rect 13527 257869 13561 257897
rect 13589 257869 13623 257897
rect 13651 257869 22437 257897
rect 22465 257869 22499 257897
rect 22527 257869 22561 257897
rect 22589 257869 22623 257897
rect 22651 257869 31437 257897
rect 31465 257869 31499 257897
rect 31527 257869 31561 257897
rect 31589 257869 31623 257897
rect 31651 257869 40437 257897
rect 40465 257869 40499 257897
rect 40527 257869 40561 257897
rect 40589 257869 40623 257897
rect 40651 257869 49437 257897
rect 49465 257869 49499 257897
rect 49527 257869 49561 257897
rect 49589 257869 49623 257897
rect 49651 257869 58437 257897
rect 58465 257869 58499 257897
rect 58527 257869 58561 257897
rect 58589 257869 58623 257897
rect 58651 257869 67437 257897
rect 67465 257869 67499 257897
rect 67527 257869 67561 257897
rect 67589 257869 67623 257897
rect 67651 257869 76437 257897
rect 76465 257869 76499 257897
rect 76527 257869 76561 257897
rect 76589 257869 76623 257897
rect 76651 257869 85437 257897
rect 85465 257869 85499 257897
rect 85527 257869 85561 257897
rect 85589 257869 85623 257897
rect 85651 257869 94437 257897
rect 94465 257869 94499 257897
rect 94527 257869 94561 257897
rect 94589 257869 94623 257897
rect 94651 257869 103437 257897
rect 103465 257869 103499 257897
rect 103527 257869 103561 257897
rect 103589 257869 103623 257897
rect 103651 257869 112437 257897
rect 112465 257869 112499 257897
rect 112527 257869 112561 257897
rect 112589 257869 112623 257897
rect 112651 257869 121437 257897
rect 121465 257869 121499 257897
rect 121527 257869 121561 257897
rect 121589 257869 121623 257897
rect 121651 257869 130437 257897
rect 130465 257869 130499 257897
rect 130527 257869 130561 257897
rect 130589 257869 130623 257897
rect 130651 257869 139437 257897
rect 139465 257869 139499 257897
rect 139527 257869 139561 257897
rect 139589 257869 139623 257897
rect 139651 257869 148437 257897
rect 148465 257869 148499 257897
rect 148527 257869 148561 257897
rect 148589 257869 148623 257897
rect 148651 257869 157437 257897
rect 157465 257869 157499 257897
rect 157527 257869 157561 257897
rect 157589 257869 157623 257897
rect 157651 257869 166437 257897
rect 166465 257869 166499 257897
rect 166527 257869 166561 257897
rect 166589 257869 166623 257897
rect 166651 257869 175437 257897
rect 175465 257869 175499 257897
rect 175527 257869 175561 257897
rect 175589 257869 175623 257897
rect 175651 257869 184437 257897
rect 184465 257869 184499 257897
rect 184527 257869 184561 257897
rect 184589 257869 184623 257897
rect 184651 257869 193437 257897
rect 193465 257869 193499 257897
rect 193527 257869 193561 257897
rect 193589 257869 193623 257897
rect 193651 257869 202437 257897
rect 202465 257869 202499 257897
rect 202527 257869 202561 257897
rect 202589 257869 202623 257897
rect 202651 257869 211437 257897
rect 211465 257869 211499 257897
rect 211527 257869 211561 257897
rect 211589 257869 211623 257897
rect 211651 257869 220437 257897
rect 220465 257869 220499 257897
rect 220527 257869 220561 257897
rect 220589 257869 220623 257897
rect 220651 257869 229437 257897
rect 229465 257869 229499 257897
rect 229527 257869 229561 257897
rect 229589 257869 229623 257897
rect 229651 257869 238437 257897
rect 238465 257869 238499 257897
rect 238527 257869 238561 257897
rect 238589 257869 238623 257897
rect 238651 257869 247437 257897
rect 247465 257869 247499 257897
rect 247527 257869 247561 257897
rect 247589 257869 247623 257897
rect 247651 257869 256437 257897
rect 256465 257869 256499 257897
rect 256527 257869 256561 257897
rect 256589 257869 256623 257897
rect 256651 257869 265437 257897
rect 265465 257869 265499 257897
rect 265527 257869 265561 257897
rect 265589 257869 265623 257897
rect 265651 257869 274437 257897
rect 274465 257869 274499 257897
rect 274527 257869 274561 257897
rect 274589 257869 274623 257897
rect 274651 257869 283437 257897
rect 283465 257869 283499 257897
rect 283527 257869 283561 257897
rect 283589 257869 283623 257897
rect 283651 257869 292437 257897
rect 292465 257869 292499 257897
rect 292527 257869 292561 257897
rect 292589 257869 292623 257897
rect 292651 257869 299736 257897
rect 299764 257869 299798 257897
rect 299826 257869 299860 257897
rect 299888 257869 299922 257897
rect 299950 257869 299998 257897
rect -6 257835 299998 257869
rect -6 257807 42 257835
rect 70 257807 104 257835
rect 132 257807 166 257835
rect 194 257807 228 257835
rect 256 257807 4437 257835
rect 4465 257807 4499 257835
rect 4527 257807 4561 257835
rect 4589 257807 4623 257835
rect 4651 257807 13437 257835
rect 13465 257807 13499 257835
rect 13527 257807 13561 257835
rect 13589 257807 13623 257835
rect 13651 257807 22437 257835
rect 22465 257807 22499 257835
rect 22527 257807 22561 257835
rect 22589 257807 22623 257835
rect 22651 257807 31437 257835
rect 31465 257807 31499 257835
rect 31527 257807 31561 257835
rect 31589 257807 31623 257835
rect 31651 257807 40437 257835
rect 40465 257807 40499 257835
rect 40527 257807 40561 257835
rect 40589 257807 40623 257835
rect 40651 257807 49437 257835
rect 49465 257807 49499 257835
rect 49527 257807 49561 257835
rect 49589 257807 49623 257835
rect 49651 257807 58437 257835
rect 58465 257807 58499 257835
rect 58527 257807 58561 257835
rect 58589 257807 58623 257835
rect 58651 257807 67437 257835
rect 67465 257807 67499 257835
rect 67527 257807 67561 257835
rect 67589 257807 67623 257835
rect 67651 257807 76437 257835
rect 76465 257807 76499 257835
rect 76527 257807 76561 257835
rect 76589 257807 76623 257835
rect 76651 257807 85437 257835
rect 85465 257807 85499 257835
rect 85527 257807 85561 257835
rect 85589 257807 85623 257835
rect 85651 257807 94437 257835
rect 94465 257807 94499 257835
rect 94527 257807 94561 257835
rect 94589 257807 94623 257835
rect 94651 257807 103437 257835
rect 103465 257807 103499 257835
rect 103527 257807 103561 257835
rect 103589 257807 103623 257835
rect 103651 257807 112437 257835
rect 112465 257807 112499 257835
rect 112527 257807 112561 257835
rect 112589 257807 112623 257835
rect 112651 257807 121437 257835
rect 121465 257807 121499 257835
rect 121527 257807 121561 257835
rect 121589 257807 121623 257835
rect 121651 257807 130437 257835
rect 130465 257807 130499 257835
rect 130527 257807 130561 257835
rect 130589 257807 130623 257835
rect 130651 257807 139437 257835
rect 139465 257807 139499 257835
rect 139527 257807 139561 257835
rect 139589 257807 139623 257835
rect 139651 257807 148437 257835
rect 148465 257807 148499 257835
rect 148527 257807 148561 257835
rect 148589 257807 148623 257835
rect 148651 257807 157437 257835
rect 157465 257807 157499 257835
rect 157527 257807 157561 257835
rect 157589 257807 157623 257835
rect 157651 257807 166437 257835
rect 166465 257807 166499 257835
rect 166527 257807 166561 257835
rect 166589 257807 166623 257835
rect 166651 257807 175437 257835
rect 175465 257807 175499 257835
rect 175527 257807 175561 257835
rect 175589 257807 175623 257835
rect 175651 257807 184437 257835
rect 184465 257807 184499 257835
rect 184527 257807 184561 257835
rect 184589 257807 184623 257835
rect 184651 257807 193437 257835
rect 193465 257807 193499 257835
rect 193527 257807 193561 257835
rect 193589 257807 193623 257835
rect 193651 257807 202437 257835
rect 202465 257807 202499 257835
rect 202527 257807 202561 257835
rect 202589 257807 202623 257835
rect 202651 257807 211437 257835
rect 211465 257807 211499 257835
rect 211527 257807 211561 257835
rect 211589 257807 211623 257835
rect 211651 257807 220437 257835
rect 220465 257807 220499 257835
rect 220527 257807 220561 257835
rect 220589 257807 220623 257835
rect 220651 257807 229437 257835
rect 229465 257807 229499 257835
rect 229527 257807 229561 257835
rect 229589 257807 229623 257835
rect 229651 257807 238437 257835
rect 238465 257807 238499 257835
rect 238527 257807 238561 257835
rect 238589 257807 238623 257835
rect 238651 257807 247437 257835
rect 247465 257807 247499 257835
rect 247527 257807 247561 257835
rect 247589 257807 247623 257835
rect 247651 257807 256437 257835
rect 256465 257807 256499 257835
rect 256527 257807 256561 257835
rect 256589 257807 256623 257835
rect 256651 257807 265437 257835
rect 265465 257807 265499 257835
rect 265527 257807 265561 257835
rect 265589 257807 265623 257835
rect 265651 257807 274437 257835
rect 274465 257807 274499 257835
rect 274527 257807 274561 257835
rect 274589 257807 274623 257835
rect 274651 257807 283437 257835
rect 283465 257807 283499 257835
rect 283527 257807 283561 257835
rect 283589 257807 283623 257835
rect 283651 257807 292437 257835
rect 292465 257807 292499 257835
rect 292527 257807 292561 257835
rect 292589 257807 292623 257835
rect 292651 257807 299736 257835
rect 299764 257807 299798 257835
rect 299826 257807 299860 257835
rect 299888 257807 299922 257835
rect 299950 257807 299998 257835
rect -6 257773 299998 257807
rect -6 257745 42 257773
rect 70 257745 104 257773
rect 132 257745 166 257773
rect 194 257745 228 257773
rect 256 257745 4437 257773
rect 4465 257745 4499 257773
rect 4527 257745 4561 257773
rect 4589 257745 4623 257773
rect 4651 257745 13437 257773
rect 13465 257745 13499 257773
rect 13527 257745 13561 257773
rect 13589 257745 13623 257773
rect 13651 257745 22437 257773
rect 22465 257745 22499 257773
rect 22527 257745 22561 257773
rect 22589 257745 22623 257773
rect 22651 257745 31437 257773
rect 31465 257745 31499 257773
rect 31527 257745 31561 257773
rect 31589 257745 31623 257773
rect 31651 257745 40437 257773
rect 40465 257745 40499 257773
rect 40527 257745 40561 257773
rect 40589 257745 40623 257773
rect 40651 257745 49437 257773
rect 49465 257745 49499 257773
rect 49527 257745 49561 257773
rect 49589 257745 49623 257773
rect 49651 257745 58437 257773
rect 58465 257745 58499 257773
rect 58527 257745 58561 257773
rect 58589 257745 58623 257773
rect 58651 257745 67437 257773
rect 67465 257745 67499 257773
rect 67527 257745 67561 257773
rect 67589 257745 67623 257773
rect 67651 257745 76437 257773
rect 76465 257745 76499 257773
rect 76527 257745 76561 257773
rect 76589 257745 76623 257773
rect 76651 257745 85437 257773
rect 85465 257745 85499 257773
rect 85527 257745 85561 257773
rect 85589 257745 85623 257773
rect 85651 257745 94437 257773
rect 94465 257745 94499 257773
rect 94527 257745 94561 257773
rect 94589 257745 94623 257773
rect 94651 257745 103437 257773
rect 103465 257745 103499 257773
rect 103527 257745 103561 257773
rect 103589 257745 103623 257773
rect 103651 257745 112437 257773
rect 112465 257745 112499 257773
rect 112527 257745 112561 257773
rect 112589 257745 112623 257773
rect 112651 257745 121437 257773
rect 121465 257745 121499 257773
rect 121527 257745 121561 257773
rect 121589 257745 121623 257773
rect 121651 257745 130437 257773
rect 130465 257745 130499 257773
rect 130527 257745 130561 257773
rect 130589 257745 130623 257773
rect 130651 257745 139437 257773
rect 139465 257745 139499 257773
rect 139527 257745 139561 257773
rect 139589 257745 139623 257773
rect 139651 257745 148437 257773
rect 148465 257745 148499 257773
rect 148527 257745 148561 257773
rect 148589 257745 148623 257773
rect 148651 257745 157437 257773
rect 157465 257745 157499 257773
rect 157527 257745 157561 257773
rect 157589 257745 157623 257773
rect 157651 257745 166437 257773
rect 166465 257745 166499 257773
rect 166527 257745 166561 257773
rect 166589 257745 166623 257773
rect 166651 257745 175437 257773
rect 175465 257745 175499 257773
rect 175527 257745 175561 257773
rect 175589 257745 175623 257773
rect 175651 257745 184437 257773
rect 184465 257745 184499 257773
rect 184527 257745 184561 257773
rect 184589 257745 184623 257773
rect 184651 257745 193437 257773
rect 193465 257745 193499 257773
rect 193527 257745 193561 257773
rect 193589 257745 193623 257773
rect 193651 257745 202437 257773
rect 202465 257745 202499 257773
rect 202527 257745 202561 257773
rect 202589 257745 202623 257773
rect 202651 257745 211437 257773
rect 211465 257745 211499 257773
rect 211527 257745 211561 257773
rect 211589 257745 211623 257773
rect 211651 257745 220437 257773
rect 220465 257745 220499 257773
rect 220527 257745 220561 257773
rect 220589 257745 220623 257773
rect 220651 257745 229437 257773
rect 229465 257745 229499 257773
rect 229527 257745 229561 257773
rect 229589 257745 229623 257773
rect 229651 257745 238437 257773
rect 238465 257745 238499 257773
rect 238527 257745 238561 257773
rect 238589 257745 238623 257773
rect 238651 257745 247437 257773
rect 247465 257745 247499 257773
rect 247527 257745 247561 257773
rect 247589 257745 247623 257773
rect 247651 257745 256437 257773
rect 256465 257745 256499 257773
rect 256527 257745 256561 257773
rect 256589 257745 256623 257773
rect 256651 257745 265437 257773
rect 265465 257745 265499 257773
rect 265527 257745 265561 257773
rect 265589 257745 265623 257773
rect 265651 257745 274437 257773
rect 274465 257745 274499 257773
rect 274527 257745 274561 257773
rect 274589 257745 274623 257773
rect 274651 257745 283437 257773
rect 283465 257745 283499 257773
rect 283527 257745 283561 257773
rect 283589 257745 283623 257773
rect 283651 257745 292437 257773
rect 292465 257745 292499 257773
rect 292527 257745 292561 257773
rect 292589 257745 292623 257773
rect 292651 257745 299736 257773
rect 299764 257745 299798 257773
rect 299826 257745 299860 257773
rect 299888 257745 299922 257773
rect 299950 257745 299998 257773
rect -6 257697 299998 257745
rect -6 254959 299998 255007
rect -6 254931 522 254959
rect 550 254931 584 254959
rect 612 254931 646 254959
rect 674 254931 708 254959
rect 736 254931 2577 254959
rect 2605 254931 2639 254959
rect 2667 254931 2701 254959
rect 2729 254931 2763 254959
rect 2791 254931 11577 254959
rect 11605 254931 11639 254959
rect 11667 254931 11701 254959
rect 11729 254931 11763 254959
rect 11791 254931 20577 254959
rect 20605 254931 20639 254959
rect 20667 254931 20701 254959
rect 20729 254931 20763 254959
rect 20791 254931 29577 254959
rect 29605 254931 29639 254959
rect 29667 254931 29701 254959
rect 29729 254931 29763 254959
rect 29791 254931 38577 254959
rect 38605 254931 38639 254959
rect 38667 254931 38701 254959
rect 38729 254931 38763 254959
rect 38791 254931 47577 254959
rect 47605 254931 47639 254959
rect 47667 254931 47701 254959
rect 47729 254931 47763 254959
rect 47791 254931 56577 254959
rect 56605 254931 56639 254959
rect 56667 254931 56701 254959
rect 56729 254931 56763 254959
rect 56791 254931 65577 254959
rect 65605 254931 65639 254959
rect 65667 254931 65701 254959
rect 65729 254931 65763 254959
rect 65791 254931 74577 254959
rect 74605 254931 74639 254959
rect 74667 254931 74701 254959
rect 74729 254931 74763 254959
rect 74791 254931 83577 254959
rect 83605 254931 83639 254959
rect 83667 254931 83701 254959
rect 83729 254931 83763 254959
rect 83791 254931 92577 254959
rect 92605 254931 92639 254959
rect 92667 254931 92701 254959
rect 92729 254931 92763 254959
rect 92791 254931 101577 254959
rect 101605 254931 101639 254959
rect 101667 254931 101701 254959
rect 101729 254931 101763 254959
rect 101791 254931 110577 254959
rect 110605 254931 110639 254959
rect 110667 254931 110701 254959
rect 110729 254931 110763 254959
rect 110791 254931 119577 254959
rect 119605 254931 119639 254959
rect 119667 254931 119701 254959
rect 119729 254931 119763 254959
rect 119791 254931 128577 254959
rect 128605 254931 128639 254959
rect 128667 254931 128701 254959
rect 128729 254931 128763 254959
rect 128791 254931 137577 254959
rect 137605 254931 137639 254959
rect 137667 254931 137701 254959
rect 137729 254931 137763 254959
rect 137791 254931 146577 254959
rect 146605 254931 146639 254959
rect 146667 254931 146701 254959
rect 146729 254931 146763 254959
rect 146791 254931 155577 254959
rect 155605 254931 155639 254959
rect 155667 254931 155701 254959
rect 155729 254931 155763 254959
rect 155791 254931 164577 254959
rect 164605 254931 164639 254959
rect 164667 254931 164701 254959
rect 164729 254931 164763 254959
rect 164791 254931 173577 254959
rect 173605 254931 173639 254959
rect 173667 254931 173701 254959
rect 173729 254931 173763 254959
rect 173791 254931 182577 254959
rect 182605 254931 182639 254959
rect 182667 254931 182701 254959
rect 182729 254931 182763 254959
rect 182791 254931 191577 254959
rect 191605 254931 191639 254959
rect 191667 254931 191701 254959
rect 191729 254931 191763 254959
rect 191791 254931 200577 254959
rect 200605 254931 200639 254959
rect 200667 254931 200701 254959
rect 200729 254931 200763 254959
rect 200791 254931 209577 254959
rect 209605 254931 209639 254959
rect 209667 254931 209701 254959
rect 209729 254931 209763 254959
rect 209791 254931 218577 254959
rect 218605 254931 218639 254959
rect 218667 254931 218701 254959
rect 218729 254931 218763 254959
rect 218791 254931 227577 254959
rect 227605 254931 227639 254959
rect 227667 254931 227701 254959
rect 227729 254931 227763 254959
rect 227791 254931 236577 254959
rect 236605 254931 236639 254959
rect 236667 254931 236701 254959
rect 236729 254931 236763 254959
rect 236791 254931 245577 254959
rect 245605 254931 245639 254959
rect 245667 254931 245701 254959
rect 245729 254931 245763 254959
rect 245791 254931 254577 254959
rect 254605 254931 254639 254959
rect 254667 254931 254701 254959
rect 254729 254931 254763 254959
rect 254791 254931 263577 254959
rect 263605 254931 263639 254959
rect 263667 254931 263701 254959
rect 263729 254931 263763 254959
rect 263791 254931 272577 254959
rect 272605 254931 272639 254959
rect 272667 254931 272701 254959
rect 272729 254931 272763 254959
rect 272791 254931 281577 254959
rect 281605 254931 281639 254959
rect 281667 254931 281701 254959
rect 281729 254931 281763 254959
rect 281791 254931 290577 254959
rect 290605 254931 290639 254959
rect 290667 254931 290701 254959
rect 290729 254931 290763 254959
rect 290791 254931 299256 254959
rect 299284 254931 299318 254959
rect 299346 254931 299380 254959
rect 299408 254931 299442 254959
rect 299470 254931 299998 254959
rect -6 254897 299998 254931
rect -6 254869 522 254897
rect 550 254869 584 254897
rect 612 254869 646 254897
rect 674 254869 708 254897
rect 736 254869 2577 254897
rect 2605 254869 2639 254897
rect 2667 254869 2701 254897
rect 2729 254869 2763 254897
rect 2791 254869 11577 254897
rect 11605 254869 11639 254897
rect 11667 254869 11701 254897
rect 11729 254869 11763 254897
rect 11791 254869 20577 254897
rect 20605 254869 20639 254897
rect 20667 254869 20701 254897
rect 20729 254869 20763 254897
rect 20791 254869 29577 254897
rect 29605 254869 29639 254897
rect 29667 254869 29701 254897
rect 29729 254869 29763 254897
rect 29791 254869 38577 254897
rect 38605 254869 38639 254897
rect 38667 254869 38701 254897
rect 38729 254869 38763 254897
rect 38791 254869 47577 254897
rect 47605 254869 47639 254897
rect 47667 254869 47701 254897
rect 47729 254869 47763 254897
rect 47791 254869 56577 254897
rect 56605 254869 56639 254897
rect 56667 254869 56701 254897
rect 56729 254869 56763 254897
rect 56791 254869 65577 254897
rect 65605 254869 65639 254897
rect 65667 254869 65701 254897
rect 65729 254869 65763 254897
rect 65791 254869 74577 254897
rect 74605 254869 74639 254897
rect 74667 254869 74701 254897
rect 74729 254869 74763 254897
rect 74791 254869 83577 254897
rect 83605 254869 83639 254897
rect 83667 254869 83701 254897
rect 83729 254869 83763 254897
rect 83791 254869 92577 254897
rect 92605 254869 92639 254897
rect 92667 254869 92701 254897
rect 92729 254869 92763 254897
rect 92791 254869 101577 254897
rect 101605 254869 101639 254897
rect 101667 254869 101701 254897
rect 101729 254869 101763 254897
rect 101791 254869 110577 254897
rect 110605 254869 110639 254897
rect 110667 254869 110701 254897
rect 110729 254869 110763 254897
rect 110791 254869 119577 254897
rect 119605 254869 119639 254897
rect 119667 254869 119701 254897
rect 119729 254869 119763 254897
rect 119791 254869 128577 254897
rect 128605 254869 128639 254897
rect 128667 254869 128701 254897
rect 128729 254869 128763 254897
rect 128791 254869 137577 254897
rect 137605 254869 137639 254897
rect 137667 254869 137701 254897
rect 137729 254869 137763 254897
rect 137791 254869 146577 254897
rect 146605 254869 146639 254897
rect 146667 254869 146701 254897
rect 146729 254869 146763 254897
rect 146791 254869 155577 254897
rect 155605 254869 155639 254897
rect 155667 254869 155701 254897
rect 155729 254869 155763 254897
rect 155791 254869 164577 254897
rect 164605 254869 164639 254897
rect 164667 254869 164701 254897
rect 164729 254869 164763 254897
rect 164791 254869 173577 254897
rect 173605 254869 173639 254897
rect 173667 254869 173701 254897
rect 173729 254869 173763 254897
rect 173791 254869 182577 254897
rect 182605 254869 182639 254897
rect 182667 254869 182701 254897
rect 182729 254869 182763 254897
rect 182791 254869 191577 254897
rect 191605 254869 191639 254897
rect 191667 254869 191701 254897
rect 191729 254869 191763 254897
rect 191791 254869 200577 254897
rect 200605 254869 200639 254897
rect 200667 254869 200701 254897
rect 200729 254869 200763 254897
rect 200791 254869 209577 254897
rect 209605 254869 209639 254897
rect 209667 254869 209701 254897
rect 209729 254869 209763 254897
rect 209791 254869 218577 254897
rect 218605 254869 218639 254897
rect 218667 254869 218701 254897
rect 218729 254869 218763 254897
rect 218791 254869 227577 254897
rect 227605 254869 227639 254897
rect 227667 254869 227701 254897
rect 227729 254869 227763 254897
rect 227791 254869 236577 254897
rect 236605 254869 236639 254897
rect 236667 254869 236701 254897
rect 236729 254869 236763 254897
rect 236791 254869 245577 254897
rect 245605 254869 245639 254897
rect 245667 254869 245701 254897
rect 245729 254869 245763 254897
rect 245791 254869 254577 254897
rect 254605 254869 254639 254897
rect 254667 254869 254701 254897
rect 254729 254869 254763 254897
rect 254791 254869 263577 254897
rect 263605 254869 263639 254897
rect 263667 254869 263701 254897
rect 263729 254869 263763 254897
rect 263791 254869 272577 254897
rect 272605 254869 272639 254897
rect 272667 254869 272701 254897
rect 272729 254869 272763 254897
rect 272791 254869 281577 254897
rect 281605 254869 281639 254897
rect 281667 254869 281701 254897
rect 281729 254869 281763 254897
rect 281791 254869 290577 254897
rect 290605 254869 290639 254897
rect 290667 254869 290701 254897
rect 290729 254869 290763 254897
rect 290791 254869 299256 254897
rect 299284 254869 299318 254897
rect 299346 254869 299380 254897
rect 299408 254869 299442 254897
rect 299470 254869 299998 254897
rect -6 254835 299998 254869
rect -6 254807 522 254835
rect 550 254807 584 254835
rect 612 254807 646 254835
rect 674 254807 708 254835
rect 736 254807 2577 254835
rect 2605 254807 2639 254835
rect 2667 254807 2701 254835
rect 2729 254807 2763 254835
rect 2791 254807 11577 254835
rect 11605 254807 11639 254835
rect 11667 254807 11701 254835
rect 11729 254807 11763 254835
rect 11791 254807 20577 254835
rect 20605 254807 20639 254835
rect 20667 254807 20701 254835
rect 20729 254807 20763 254835
rect 20791 254807 29577 254835
rect 29605 254807 29639 254835
rect 29667 254807 29701 254835
rect 29729 254807 29763 254835
rect 29791 254807 38577 254835
rect 38605 254807 38639 254835
rect 38667 254807 38701 254835
rect 38729 254807 38763 254835
rect 38791 254807 47577 254835
rect 47605 254807 47639 254835
rect 47667 254807 47701 254835
rect 47729 254807 47763 254835
rect 47791 254807 56577 254835
rect 56605 254807 56639 254835
rect 56667 254807 56701 254835
rect 56729 254807 56763 254835
rect 56791 254807 65577 254835
rect 65605 254807 65639 254835
rect 65667 254807 65701 254835
rect 65729 254807 65763 254835
rect 65791 254807 74577 254835
rect 74605 254807 74639 254835
rect 74667 254807 74701 254835
rect 74729 254807 74763 254835
rect 74791 254807 83577 254835
rect 83605 254807 83639 254835
rect 83667 254807 83701 254835
rect 83729 254807 83763 254835
rect 83791 254807 92577 254835
rect 92605 254807 92639 254835
rect 92667 254807 92701 254835
rect 92729 254807 92763 254835
rect 92791 254807 101577 254835
rect 101605 254807 101639 254835
rect 101667 254807 101701 254835
rect 101729 254807 101763 254835
rect 101791 254807 110577 254835
rect 110605 254807 110639 254835
rect 110667 254807 110701 254835
rect 110729 254807 110763 254835
rect 110791 254807 119577 254835
rect 119605 254807 119639 254835
rect 119667 254807 119701 254835
rect 119729 254807 119763 254835
rect 119791 254807 128577 254835
rect 128605 254807 128639 254835
rect 128667 254807 128701 254835
rect 128729 254807 128763 254835
rect 128791 254807 137577 254835
rect 137605 254807 137639 254835
rect 137667 254807 137701 254835
rect 137729 254807 137763 254835
rect 137791 254807 146577 254835
rect 146605 254807 146639 254835
rect 146667 254807 146701 254835
rect 146729 254807 146763 254835
rect 146791 254807 155577 254835
rect 155605 254807 155639 254835
rect 155667 254807 155701 254835
rect 155729 254807 155763 254835
rect 155791 254807 164577 254835
rect 164605 254807 164639 254835
rect 164667 254807 164701 254835
rect 164729 254807 164763 254835
rect 164791 254807 173577 254835
rect 173605 254807 173639 254835
rect 173667 254807 173701 254835
rect 173729 254807 173763 254835
rect 173791 254807 182577 254835
rect 182605 254807 182639 254835
rect 182667 254807 182701 254835
rect 182729 254807 182763 254835
rect 182791 254807 191577 254835
rect 191605 254807 191639 254835
rect 191667 254807 191701 254835
rect 191729 254807 191763 254835
rect 191791 254807 200577 254835
rect 200605 254807 200639 254835
rect 200667 254807 200701 254835
rect 200729 254807 200763 254835
rect 200791 254807 209577 254835
rect 209605 254807 209639 254835
rect 209667 254807 209701 254835
rect 209729 254807 209763 254835
rect 209791 254807 218577 254835
rect 218605 254807 218639 254835
rect 218667 254807 218701 254835
rect 218729 254807 218763 254835
rect 218791 254807 227577 254835
rect 227605 254807 227639 254835
rect 227667 254807 227701 254835
rect 227729 254807 227763 254835
rect 227791 254807 236577 254835
rect 236605 254807 236639 254835
rect 236667 254807 236701 254835
rect 236729 254807 236763 254835
rect 236791 254807 245577 254835
rect 245605 254807 245639 254835
rect 245667 254807 245701 254835
rect 245729 254807 245763 254835
rect 245791 254807 254577 254835
rect 254605 254807 254639 254835
rect 254667 254807 254701 254835
rect 254729 254807 254763 254835
rect 254791 254807 263577 254835
rect 263605 254807 263639 254835
rect 263667 254807 263701 254835
rect 263729 254807 263763 254835
rect 263791 254807 272577 254835
rect 272605 254807 272639 254835
rect 272667 254807 272701 254835
rect 272729 254807 272763 254835
rect 272791 254807 281577 254835
rect 281605 254807 281639 254835
rect 281667 254807 281701 254835
rect 281729 254807 281763 254835
rect 281791 254807 290577 254835
rect 290605 254807 290639 254835
rect 290667 254807 290701 254835
rect 290729 254807 290763 254835
rect 290791 254807 299256 254835
rect 299284 254807 299318 254835
rect 299346 254807 299380 254835
rect 299408 254807 299442 254835
rect 299470 254807 299998 254835
rect -6 254773 299998 254807
rect -6 254745 522 254773
rect 550 254745 584 254773
rect 612 254745 646 254773
rect 674 254745 708 254773
rect 736 254745 2577 254773
rect 2605 254745 2639 254773
rect 2667 254745 2701 254773
rect 2729 254745 2763 254773
rect 2791 254745 11577 254773
rect 11605 254745 11639 254773
rect 11667 254745 11701 254773
rect 11729 254745 11763 254773
rect 11791 254745 20577 254773
rect 20605 254745 20639 254773
rect 20667 254745 20701 254773
rect 20729 254745 20763 254773
rect 20791 254745 29577 254773
rect 29605 254745 29639 254773
rect 29667 254745 29701 254773
rect 29729 254745 29763 254773
rect 29791 254745 38577 254773
rect 38605 254745 38639 254773
rect 38667 254745 38701 254773
rect 38729 254745 38763 254773
rect 38791 254745 47577 254773
rect 47605 254745 47639 254773
rect 47667 254745 47701 254773
rect 47729 254745 47763 254773
rect 47791 254745 56577 254773
rect 56605 254745 56639 254773
rect 56667 254745 56701 254773
rect 56729 254745 56763 254773
rect 56791 254745 65577 254773
rect 65605 254745 65639 254773
rect 65667 254745 65701 254773
rect 65729 254745 65763 254773
rect 65791 254745 74577 254773
rect 74605 254745 74639 254773
rect 74667 254745 74701 254773
rect 74729 254745 74763 254773
rect 74791 254745 83577 254773
rect 83605 254745 83639 254773
rect 83667 254745 83701 254773
rect 83729 254745 83763 254773
rect 83791 254745 92577 254773
rect 92605 254745 92639 254773
rect 92667 254745 92701 254773
rect 92729 254745 92763 254773
rect 92791 254745 101577 254773
rect 101605 254745 101639 254773
rect 101667 254745 101701 254773
rect 101729 254745 101763 254773
rect 101791 254745 110577 254773
rect 110605 254745 110639 254773
rect 110667 254745 110701 254773
rect 110729 254745 110763 254773
rect 110791 254745 119577 254773
rect 119605 254745 119639 254773
rect 119667 254745 119701 254773
rect 119729 254745 119763 254773
rect 119791 254745 128577 254773
rect 128605 254745 128639 254773
rect 128667 254745 128701 254773
rect 128729 254745 128763 254773
rect 128791 254745 137577 254773
rect 137605 254745 137639 254773
rect 137667 254745 137701 254773
rect 137729 254745 137763 254773
rect 137791 254745 146577 254773
rect 146605 254745 146639 254773
rect 146667 254745 146701 254773
rect 146729 254745 146763 254773
rect 146791 254745 155577 254773
rect 155605 254745 155639 254773
rect 155667 254745 155701 254773
rect 155729 254745 155763 254773
rect 155791 254745 164577 254773
rect 164605 254745 164639 254773
rect 164667 254745 164701 254773
rect 164729 254745 164763 254773
rect 164791 254745 173577 254773
rect 173605 254745 173639 254773
rect 173667 254745 173701 254773
rect 173729 254745 173763 254773
rect 173791 254745 182577 254773
rect 182605 254745 182639 254773
rect 182667 254745 182701 254773
rect 182729 254745 182763 254773
rect 182791 254745 191577 254773
rect 191605 254745 191639 254773
rect 191667 254745 191701 254773
rect 191729 254745 191763 254773
rect 191791 254745 200577 254773
rect 200605 254745 200639 254773
rect 200667 254745 200701 254773
rect 200729 254745 200763 254773
rect 200791 254745 209577 254773
rect 209605 254745 209639 254773
rect 209667 254745 209701 254773
rect 209729 254745 209763 254773
rect 209791 254745 218577 254773
rect 218605 254745 218639 254773
rect 218667 254745 218701 254773
rect 218729 254745 218763 254773
rect 218791 254745 227577 254773
rect 227605 254745 227639 254773
rect 227667 254745 227701 254773
rect 227729 254745 227763 254773
rect 227791 254745 236577 254773
rect 236605 254745 236639 254773
rect 236667 254745 236701 254773
rect 236729 254745 236763 254773
rect 236791 254745 245577 254773
rect 245605 254745 245639 254773
rect 245667 254745 245701 254773
rect 245729 254745 245763 254773
rect 245791 254745 254577 254773
rect 254605 254745 254639 254773
rect 254667 254745 254701 254773
rect 254729 254745 254763 254773
rect 254791 254745 263577 254773
rect 263605 254745 263639 254773
rect 263667 254745 263701 254773
rect 263729 254745 263763 254773
rect 263791 254745 272577 254773
rect 272605 254745 272639 254773
rect 272667 254745 272701 254773
rect 272729 254745 272763 254773
rect 272791 254745 281577 254773
rect 281605 254745 281639 254773
rect 281667 254745 281701 254773
rect 281729 254745 281763 254773
rect 281791 254745 290577 254773
rect 290605 254745 290639 254773
rect 290667 254745 290701 254773
rect 290729 254745 290763 254773
rect 290791 254745 299256 254773
rect 299284 254745 299318 254773
rect 299346 254745 299380 254773
rect 299408 254745 299442 254773
rect 299470 254745 299998 254773
rect -6 254697 299998 254745
rect -6 248959 299998 249007
rect -6 248931 42 248959
rect 70 248931 104 248959
rect 132 248931 166 248959
rect 194 248931 228 248959
rect 256 248931 4437 248959
rect 4465 248931 4499 248959
rect 4527 248931 4561 248959
rect 4589 248931 4623 248959
rect 4651 248931 13437 248959
rect 13465 248931 13499 248959
rect 13527 248931 13561 248959
rect 13589 248931 13623 248959
rect 13651 248931 22437 248959
rect 22465 248931 22499 248959
rect 22527 248931 22561 248959
rect 22589 248931 22623 248959
rect 22651 248931 24939 248959
rect 24967 248931 25001 248959
rect 25029 248931 31437 248959
rect 31465 248931 31499 248959
rect 31527 248931 31561 248959
rect 31589 248931 31623 248959
rect 31651 248931 40299 248959
rect 40327 248931 40361 248959
rect 40389 248931 55659 248959
rect 55687 248931 55721 248959
rect 55749 248931 71019 248959
rect 71047 248931 71081 248959
rect 71109 248931 86379 248959
rect 86407 248931 86441 248959
rect 86469 248931 101739 248959
rect 101767 248931 101801 248959
rect 101829 248931 117099 248959
rect 117127 248931 117161 248959
rect 117189 248931 132459 248959
rect 132487 248931 132521 248959
rect 132549 248931 147819 248959
rect 147847 248931 147881 248959
rect 147909 248931 163179 248959
rect 163207 248931 163241 248959
rect 163269 248931 178539 248959
rect 178567 248931 178601 248959
rect 178629 248931 193899 248959
rect 193927 248931 193961 248959
rect 193989 248931 209259 248959
rect 209287 248931 209321 248959
rect 209349 248931 224619 248959
rect 224647 248931 224681 248959
rect 224709 248931 239979 248959
rect 240007 248931 240041 248959
rect 240069 248931 256437 248959
rect 256465 248931 256499 248959
rect 256527 248931 256561 248959
rect 256589 248931 256623 248959
rect 256651 248931 265437 248959
rect 265465 248931 265499 248959
rect 265527 248931 265561 248959
rect 265589 248931 265623 248959
rect 265651 248931 274437 248959
rect 274465 248931 274499 248959
rect 274527 248931 274561 248959
rect 274589 248931 274623 248959
rect 274651 248931 283437 248959
rect 283465 248931 283499 248959
rect 283527 248931 283561 248959
rect 283589 248931 283623 248959
rect 283651 248931 292437 248959
rect 292465 248931 292499 248959
rect 292527 248931 292561 248959
rect 292589 248931 292623 248959
rect 292651 248931 299736 248959
rect 299764 248931 299798 248959
rect 299826 248931 299860 248959
rect 299888 248931 299922 248959
rect 299950 248931 299998 248959
rect -6 248897 299998 248931
rect -6 248869 42 248897
rect 70 248869 104 248897
rect 132 248869 166 248897
rect 194 248869 228 248897
rect 256 248869 4437 248897
rect 4465 248869 4499 248897
rect 4527 248869 4561 248897
rect 4589 248869 4623 248897
rect 4651 248869 13437 248897
rect 13465 248869 13499 248897
rect 13527 248869 13561 248897
rect 13589 248869 13623 248897
rect 13651 248869 22437 248897
rect 22465 248869 22499 248897
rect 22527 248869 22561 248897
rect 22589 248869 22623 248897
rect 22651 248869 24939 248897
rect 24967 248869 25001 248897
rect 25029 248869 31437 248897
rect 31465 248869 31499 248897
rect 31527 248869 31561 248897
rect 31589 248869 31623 248897
rect 31651 248869 40299 248897
rect 40327 248869 40361 248897
rect 40389 248869 55659 248897
rect 55687 248869 55721 248897
rect 55749 248869 71019 248897
rect 71047 248869 71081 248897
rect 71109 248869 86379 248897
rect 86407 248869 86441 248897
rect 86469 248869 101739 248897
rect 101767 248869 101801 248897
rect 101829 248869 117099 248897
rect 117127 248869 117161 248897
rect 117189 248869 132459 248897
rect 132487 248869 132521 248897
rect 132549 248869 147819 248897
rect 147847 248869 147881 248897
rect 147909 248869 163179 248897
rect 163207 248869 163241 248897
rect 163269 248869 178539 248897
rect 178567 248869 178601 248897
rect 178629 248869 193899 248897
rect 193927 248869 193961 248897
rect 193989 248869 209259 248897
rect 209287 248869 209321 248897
rect 209349 248869 224619 248897
rect 224647 248869 224681 248897
rect 224709 248869 239979 248897
rect 240007 248869 240041 248897
rect 240069 248869 256437 248897
rect 256465 248869 256499 248897
rect 256527 248869 256561 248897
rect 256589 248869 256623 248897
rect 256651 248869 265437 248897
rect 265465 248869 265499 248897
rect 265527 248869 265561 248897
rect 265589 248869 265623 248897
rect 265651 248869 274437 248897
rect 274465 248869 274499 248897
rect 274527 248869 274561 248897
rect 274589 248869 274623 248897
rect 274651 248869 283437 248897
rect 283465 248869 283499 248897
rect 283527 248869 283561 248897
rect 283589 248869 283623 248897
rect 283651 248869 292437 248897
rect 292465 248869 292499 248897
rect 292527 248869 292561 248897
rect 292589 248869 292623 248897
rect 292651 248869 299736 248897
rect 299764 248869 299798 248897
rect 299826 248869 299860 248897
rect 299888 248869 299922 248897
rect 299950 248869 299998 248897
rect -6 248835 299998 248869
rect -6 248807 42 248835
rect 70 248807 104 248835
rect 132 248807 166 248835
rect 194 248807 228 248835
rect 256 248807 4437 248835
rect 4465 248807 4499 248835
rect 4527 248807 4561 248835
rect 4589 248807 4623 248835
rect 4651 248807 13437 248835
rect 13465 248807 13499 248835
rect 13527 248807 13561 248835
rect 13589 248807 13623 248835
rect 13651 248807 22437 248835
rect 22465 248807 22499 248835
rect 22527 248807 22561 248835
rect 22589 248807 22623 248835
rect 22651 248807 24939 248835
rect 24967 248807 25001 248835
rect 25029 248807 31437 248835
rect 31465 248807 31499 248835
rect 31527 248807 31561 248835
rect 31589 248807 31623 248835
rect 31651 248807 40299 248835
rect 40327 248807 40361 248835
rect 40389 248807 55659 248835
rect 55687 248807 55721 248835
rect 55749 248807 71019 248835
rect 71047 248807 71081 248835
rect 71109 248807 86379 248835
rect 86407 248807 86441 248835
rect 86469 248807 101739 248835
rect 101767 248807 101801 248835
rect 101829 248807 117099 248835
rect 117127 248807 117161 248835
rect 117189 248807 132459 248835
rect 132487 248807 132521 248835
rect 132549 248807 147819 248835
rect 147847 248807 147881 248835
rect 147909 248807 163179 248835
rect 163207 248807 163241 248835
rect 163269 248807 178539 248835
rect 178567 248807 178601 248835
rect 178629 248807 193899 248835
rect 193927 248807 193961 248835
rect 193989 248807 209259 248835
rect 209287 248807 209321 248835
rect 209349 248807 224619 248835
rect 224647 248807 224681 248835
rect 224709 248807 239979 248835
rect 240007 248807 240041 248835
rect 240069 248807 256437 248835
rect 256465 248807 256499 248835
rect 256527 248807 256561 248835
rect 256589 248807 256623 248835
rect 256651 248807 265437 248835
rect 265465 248807 265499 248835
rect 265527 248807 265561 248835
rect 265589 248807 265623 248835
rect 265651 248807 274437 248835
rect 274465 248807 274499 248835
rect 274527 248807 274561 248835
rect 274589 248807 274623 248835
rect 274651 248807 283437 248835
rect 283465 248807 283499 248835
rect 283527 248807 283561 248835
rect 283589 248807 283623 248835
rect 283651 248807 292437 248835
rect 292465 248807 292499 248835
rect 292527 248807 292561 248835
rect 292589 248807 292623 248835
rect 292651 248807 299736 248835
rect 299764 248807 299798 248835
rect 299826 248807 299860 248835
rect 299888 248807 299922 248835
rect 299950 248807 299998 248835
rect -6 248773 299998 248807
rect -6 248745 42 248773
rect 70 248745 104 248773
rect 132 248745 166 248773
rect 194 248745 228 248773
rect 256 248745 4437 248773
rect 4465 248745 4499 248773
rect 4527 248745 4561 248773
rect 4589 248745 4623 248773
rect 4651 248745 13437 248773
rect 13465 248745 13499 248773
rect 13527 248745 13561 248773
rect 13589 248745 13623 248773
rect 13651 248745 22437 248773
rect 22465 248745 22499 248773
rect 22527 248745 22561 248773
rect 22589 248745 22623 248773
rect 22651 248745 24939 248773
rect 24967 248745 25001 248773
rect 25029 248745 31437 248773
rect 31465 248745 31499 248773
rect 31527 248745 31561 248773
rect 31589 248745 31623 248773
rect 31651 248745 40299 248773
rect 40327 248745 40361 248773
rect 40389 248745 55659 248773
rect 55687 248745 55721 248773
rect 55749 248745 71019 248773
rect 71047 248745 71081 248773
rect 71109 248745 86379 248773
rect 86407 248745 86441 248773
rect 86469 248745 101739 248773
rect 101767 248745 101801 248773
rect 101829 248745 117099 248773
rect 117127 248745 117161 248773
rect 117189 248745 132459 248773
rect 132487 248745 132521 248773
rect 132549 248745 147819 248773
rect 147847 248745 147881 248773
rect 147909 248745 163179 248773
rect 163207 248745 163241 248773
rect 163269 248745 178539 248773
rect 178567 248745 178601 248773
rect 178629 248745 193899 248773
rect 193927 248745 193961 248773
rect 193989 248745 209259 248773
rect 209287 248745 209321 248773
rect 209349 248745 224619 248773
rect 224647 248745 224681 248773
rect 224709 248745 239979 248773
rect 240007 248745 240041 248773
rect 240069 248745 256437 248773
rect 256465 248745 256499 248773
rect 256527 248745 256561 248773
rect 256589 248745 256623 248773
rect 256651 248745 265437 248773
rect 265465 248745 265499 248773
rect 265527 248745 265561 248773
rect 265589 248745 265623 248773
rect 265651 248745 274437 248773
rect 274465 248745 274499 248773
rect 274527 248745 274561 248773
rect 274589 248745 274623 248773
rect 274651 248745 283437 248773
rect 283465 248745 283499 248773
rect 283527 248745 283561 248773
rect 283589 248745 283623 248773
rect 283651 248745 292437 248773
rect 292465 248745 292499 248773
rect 292527 248745 292561 248773
rect 292589 248745 292623 248773
rect 292651 248745 299736 248773
rect 299764 248745 299798 248773
rect 299826 248745 299860 248773
rect 299888 248745 299922 248773
rect 299950 248745 299998 248773
rect -6 248697 299998 248745
rect -6 245959 299998 246007
rect -6 245931 522 245959
rect 550 245931 584 245959
rect 612 245931 646 245959
rect 674 245931 708 245959
rect 736 245931 2577 245959
rect 2605 245931 2639 245959
rect 2667 245931 2701 245959
rect 2729 245931 2763 245959
rect 2791 245931 11577 245959
rect 11605 245931 11639 245959
rect 11667 245931 11701 245959
rect 11729 245931 11763 245959
rect 11791 245931 17259 245959
rect 17287 245931 17321 245959
rect 17349 245931 20577 245959
rect 20605 245931 20639 245959
rect 20667 245931 20701 245959
rect 20729 245931 20763 245959
rect 20791 245931 29577 245959
rect 29605 245931 29639 245959
rect 29667 245931 29701 245959
rect 29729 245931 29763 245959
rect 29791 245931 32619 245959
rect 32647 245931 32681 245959
rect 32709 245931 47979 245959
rect 48007 245931 48041 245959
rect 48069 245931 63339 245959
rect 63367 245931 63401 245959
rect 63429 245931 78699 245959
rect 78727 245931 78761 245959
rect 78789 245931 94059 245959
rect 94087 245931 94121 245959
rect 94149 245931 109419 245959
rect 109447 245931 109481 245959
rect 109509 245931 124779 245959
rect 124807 245931 124841 245959
rect 124869 245931 140139 245959
rect 140167 245931 140201 245959
rect 140229 245931 155499 245959
rect 155527 245931 155561 245959
rect 155589 245931 170859 245959
rect 170887 245931 170921 245959
rect 170949 245931 186219 245959
rect 186247 245931 186281 245959
rect 186309 245931 201579 245959
rect 201607 245931 201641 245959
rect 201669 245931 216939 245959
rect 216967 245931 217001 245959
rect 217029 245931 232299 245959
rect 232327 245931 232361 245959
rect 232389 245931 247659 245959
rect 247687 245931 247721 245959
rect 247749 245931 254577 245959
rect 254605 245931 254639 245959
rect 254667 245931 254701 245959
rect 254729 245931 254763 245959
rect 254791 245931 263577 245959
rect 263605 245931 263639 245959
rect 263667 245931 263701 245959
rect 263729 245931 263763 245959
rect 263791 245931 272577 245959
rect 272605 245931 272639 245959
rect 272667 245931 272701 245959
rect 272729 245931 272763 245959
rect 272791 245931 281577 245959
rect 281605 245931 281639 245959
rect 281667 245931 281701 245959
rect 281729 245931 281763 245959
rect 281791 245931 290577 245959
rect 290605 245931 290639 245959
rect 290667 245931 290701 245959
rect 290729 245931 290763 245959
rect 290791 245931 299256 245959
rect 299284 245931 299318 245959
rect 299346 245931 299380 245959
rect 299408 245931 299442 245959
rect 299470 245931 299998 245959
rect -6 245897 299998 245931
rect -6 245869 522 245897
rect 550 245869 584 245897
rect 612 245869 646 245897
rect 674 245869 708 245897
rect 736 245869 2577 245897
rect 2605 245869 2639 245897
rect 2667 245869 2701 245897
rect 2729 245869 2763 245897
rect 2791 245869 11577 245897
rect 11605 245869 11639 245897
rect 11667 245869 11701 245897
rect 11729 245869 11763 245897
rect 11791 245869 17259 245897
rect 17287 245869 17321 245897
rect 17349 245869 20577 245897
rect 20605 245869 20639 245897
rect 20667 245869 20701 245897
rect 20729 245869 20763 245897
rect 20791 245869 29577 245897
rect 29605 245869 29639 245897
rect 29667 245869 29701 245897
rect 29729 245869 29763 245897
rect 29791 245869 32619 245897
rect 32647 245869 32681 245897
rect 32709 245869 47979 245897
rect 48007 245869 48041 245897
rect 48069 245869 63339 245897
rect 63367 245869 63401 245897
rect 63429 245869 78699 245897
rect 78727 245869 78761 245897
rect 78789 245869 94059 245897
rect 94087 245869 94121 245897
rect 94149 245869 109419 245897
rect 109447 245869 109481 245897
rect 109509 245869 124779 245897
rect 124807 245869 124841 245897
rect 124869 245869 140139 245897
rect 140167 245869 140201 245897
rect 140229 245869 155499 245897
rect 155527 245869 155561 245897
rect 155589 245869 170859 245897
rect 170887 245869 170921 245897
rect 170949 245869 186219 245897
rect 186247 245869 186281 245897
rect 186309 245869 201579 245897
rect 201607 245869 201641 245897
rect 201669 245869 216939 245897
rect 216967 245869 217001 245897
rect 217029 245869 232299 245897
rect 232327 245869 232361 245897
rect 232389 245869 247659 245897
rect 247687 245869 247721 245897
rect 247749 245869 254577 245897
rect 254605 245869 254639 245897
rect 254667 245869 254701 245897
rect 254729 245869 254763 245897
rect 254791 245869 263577 245897
rect 263605 245869 263639 245897
rect 263667 245869 263701 245897
rect 263729 245869 263763 245897
rect 263791 245869 272577 245897
rect 272605 245869 272639 245897
rect 272667 245869 272701 245897
rect 272729 245869 272763 245897
rect 272791 245869 281577 245897
rect 281605 245869 281639 245897
rect 281667 245869 281701 245897
rect 281729 245869 281763 245897
rect 281791 245869 290577 245897
rect 290605 245869 290639 245897
rect 290667 245869 290701 245897
rect 290729 245869 290763 245897
rect 290791 245869 299256 245897
rect 299284 245869 299318 245897
rect 299346 245869 299380 245897
rect 299408 245869 299442 245897
rect 299470 245869 299998 245897
rect -6 245835 299998 245869
rect -6 245807 522 245835
rect 550 245807 584 245835
rect 612 245807 646 245835
rect 674 245807 708 245835
rect 736 245807 2577 245835
rect 2605 245807 2639 245835
rect 2667 245807 2701 245835
rect 2729 245807 2763 245835
rect 2791 245807 11577 245835
rect 11605 245807 11639 245835
rect 11667 245807 11701 245835
rect 11729 245807 11763 245835
rect 11791 245807 17259 245835
rect 17287 245807 17321 245835
rect 17349 245807 20577 245835
rect 20605 245807 20639 245835
rect 20667 245807 20701 245835
rect 20729 245807 20763 245835
rect 20791 245807 29577 245835
rect 29605 245807 29639 245835
rect 29667 245807 29701 245835
rect 29729 245807 29763 245835
rect 29791 245807 32619 245835
rect 32647 245807 32681 245835
rect 32709 245807 47979 245835
rect 48007 245807 48041 245835
rect 48069 245807 63339 245835
rect 63367 245807 63401 245835
rect 63429 245807 78699 245835
rect 78727 245807 78761 245835
rect 78789 245807 94059 245835
rect 94087 245807 94121 245835
rect 94149 245807 109419 245835
rect 109447 245807 109481 245835
rect 109509 245807 124779 245835
rect 124807 245807 124841 245835
rect 124869 245807 140139 245835
rect 140167 245807 140201 245835
rect 140229 245807 155499 245835
rect 155527 245807 155561 245835
rect 155589 245807 170859 245835
rect 170887 245807 170921 245835
rect 170949 245807 186219 245835
rect 186247 245807 186281 245835
rect 186309 245807 201579 245835
rect 201607 245807 201641 245835
rect 201669 245807 216939 245835
rect 216967 245807 217001 245835
rect 217029 245807 232299 245835
rect 232327 245807 232361 245835
rect 232389 245807 247659 245835
rect 247687 245807 247721 245835
rect 247749 245807 254577 245835
rect 254605 245807 254639 245835
rect 254667 245807 254701 245835
rect 254729 245807 254763 245835
rect 254791 245807 263577 245835
rect 263605 245807 263639 245835
rect 263667 245807 263701 245835
rect 263729 245807 263763 245835
rect 263791 245807 272577 245835
rect 272605 245807 272639 245835
rect 272667 245807 272701 245835
rect 272729 245807 272763 245835
rect 272791 245807 281577 245835
rect 281605 245807 281639 245835
rect 281667 245807 281701 245835
rect 281729 245807 281763 245835
rect 281791 245807 290577 245835
rect 290605 245807 290639 245835
rect 290667 245807 290701 245835
rect 290729 245807 290763 245835
rect 290791 245807 299256 245835
rect 299284 245807 299318 245835
rect 299346 245807 299380 245835
rect 299408 245807 299442 245835
rect 299470 245807 299998 245835
rect -6 245773 299998 245807
rect -6 245745 522 245773
rect 550 245745 584 245773
rect 612 245745 646 245773
rect 674 245745 708 245773
rect 736 245745 2577 245773
rect 2605 245745 2639 245773
rect 2667 245745 2701 245773
rect 2729 245745 2763 245773
rect 2791 245745 11577 245773
rect 11605 245745 11639 245773
rect 11667 245745 11701 245773
rect 11729 245745 11763 245773
rect 11791 245745 17259 245773
rect 17287 245745 17321 245773
rect 17349 245745 20577 245773
rect 20605 245745 20639 245773
rect 20667 245745 20701 245773
rect 20729 245745 20763 245773
rect 20791 245745 29577 245773
rect 29605 245745 29639 245773
rect 29667 245745 29701 245773
rect 29729 245745 29763 245773
rect 29791 245745 32619 245773
rect 32647 245745 32681 245773
rect 32709 245745 47979 245773
rect 48007 245745 48041 245773
rect 48069 245745 63339 245773
rect 63367 245745 63401 245773
rect 63429 245745 78699 245773
rect 78727 245745 78761 245773
rect 78789 245745 94059 245773
rect 94087 245745 94121 245773
rect 94149 245745 109419 245773
rect 109447 245745 109481 245773
rect 109509 245745 124779 245773
rect 124807 245745 124841 245773
rect 124869 245745 140139 245773
rect 140167 245745 140201 245773
rect 140229 245745 155499 245773
rect 155527 245745 155561 245773
rect 155589 245745 170859 245773
rect 170887 245745 170921 245773
rect 170949 245745 186219 245773
rect 186247 245745 186281 245773
rect 186309 245745 201579 245773
rect 201607 245745 201641 245773
rect 201669 245745 216939 245773
rect 216967 245745 217001 245773
rect 217029 245745 232299 245773
rect 232327 245745 232361 245773
rect 232389 245745 247659 245773
rect 247687 245745 247721 245773
rect 247749 245745 254577 245773
rect 254605 245745 254639 245773
rect 254667 245745 254701 245773
rect 254729 245745 254763 245773
rect 254791 245745 263577 245773
rect 263605 245745 263639 245773
rect 263667 245745 263701 245773
rect 263729 245745 263763 245773
rect 263791 245745 272577 245773
rect 272605 245745 272639 245773
rect 272667 245745 272701 245773
rect 272729 245745 272763 245773
rect 272791 245745 281577 245773
rect 281605 245745 281639 245773
rect 281667 245745 281701 245773
rect 281729 245745 281763 245773
rect 281791 245745 290577 245773
rect 290605 245745 290639 245773
rect 290667 245745 290701 245773
rect 290729 245745 290763 245773
rect 290791 245745 299256 245773
rect 299284 245745 299318 245773
rect 299346 245745 299380 245773
rect 299408 245745 299442 245773
rect 299470 245745 299998 245773
rect -6 245697 299998 245745
rect -6 239959 299998 240007
rect -6 239931 42 239959
rect 70 239931 104 239959
rect 132 239931 166 239959
rect 194 239931 228 239959
rect 256 239931 4437 239959
rect 4465 239931 4499 239959
rect 4527 239931 4561 239959
rect 4589 239931 4623 239959
rect 4651 239931 13437 239959
rect 13465 239931 13499 239959
rect 13527 239931 13561 239959
rect 13589 239931 13623 239959
rect 13651 239931 22437 239959
rect 22465 239931 22499 239959
rect 22527 239931 22561 239959
rect 22589 239931 22623 239959
rect 22651 239931 24939 239959
rect 24967 239931 25001 239959
rect 25029 239931 31437 239959
rect 31465 239931 31499 239959
rect 31527 239931 31561 239959
rect 31589 239931 31623 239959
rect 31651 239931 40299 239959
rect 40327 239931 40361 239959
rect 40389 239931 55659 239959
rect 55687 239931 55721 239959
rect 55749 239931 71019 239959
rect 71047 239931 71081 239959
rect 71109 239931 86379 239959
rect 86407 239931 86441 239959
rect 86469 239931 101739 239959
rect 101767 239931 101801 239959
rect 101829 239931 117099 239959
rect 117127 239931 117161 239959
rect 117189 239931 132459 239959
rect 132487 239931 132521 239959
rect 132549 239931 147819 239959
rect 147847 239931 147881 239959
rect 147909 239931 163179 239959
rect 163207 239931 163241 239959
rect 163269 239931 178539 239959
rect 178567 239931 178601 239959
rect 178629 239931 193899 239959
rect 193927 239931 193961 239959
rect 193989 239931 209259 239959
rect 209287 239931 209321 239959
rect 209349 239931 224619 239959
rect 224647 239931 224681 239959
rect 224709 239931 239979 239959
rect 240007 239931 240041 239959
rect 240069 239931 256437 239959
rect 256465 239931 256499 239959
rect 256527 239931 256561 239959
rect 256589 239931 256623 239959
rect 256651 239931 265437 239959
rect 265465 239931 265499 239959
rect 265527 239931 265561 239959
rect 265589 239931 265623 239959
rect 265651 239931 274437 239959
rect 274465 239931 274499 239959
rect 274527 239931 274561 239959
rect 274589 239931 274623 239959
rect 274651 239931 283437 239959
rect 283465 239931 283499 239959
rect 283527 239931 283561 239959
rect 283589 239931 283623 239959
rect 283651 239931 292437 239959
rect 292465 239931 292499 239959
rect 292527 239931 292561 239959
rect 292589 239931 292623 239959
rect 292651 239931 299736 239959
rect 299764 239931 299798 239959
rect 299826 239931 299860 239959
rect 299888 239931 299922 239959
rect 299950 239931 299998 239959
rect -6 239897 299998 239931
rect -6 239869 42 239897
rect 70 239869 104 239897
rect 132 239869 166 239897
rect 194 239869 228 239897
rect 256 239869 4437 239897
rect 4465 239869 4499 239897
rect 4527 239869 4561 239897
rect 4589 239869 4623 239897
rect 4651 239869 13437 239897
rect 13465 239869 13499 239897
rect 13527 239869 13561 239897
rect 13589 239869 13623 239897
rect 13651 239869 22437 239897
rect 22465 239869 22499 239897
rect 22527 239869 22561 239897
rect 22589 239869 22623 239897
rect 22651 239869 24939 239897
rect 24967 239869 25001 239897
rect 25029 239869 31437 239897
rect 31465 239869 31499 239897
rect 31527 239869 31561 239897
rect 31589 239869 31623 239897
rect 31651 239869 40299 239897
rect 40327 239869 40361 239897
rect 40389 239869 55659 239897
rect 55687 239869 55721 239897
rect 55749 239869 71019 239897
rect 71047 239869 71081 239897
rect 71109 239869 86379 239897
rect 86407 239869 86441 239897
rect 86469 239869 101739 239897
rect 101767 239869 101801 239897
rect 101829 239869 117099 239897
rect 117127 239869 117161 239897
rect 117189 239869 132459 239897
rect 132487 239869 132521 239897
rect 132549 239869 147819 239897
rect 147847 239869 147881 239897
rect 147909 239869 163179 239897
rect 163207 239869 163241 239897
rect 163269 239869 178539 239897
rect 178567 239869 178601 239897
rect 178629 239869 193899 239897
rect 193927 239869 193961 239897
rect 193989 239869 209259 239897
rect 209287 239869 209321 239897
rect 209349 239869 224619 239897
rect 224647 239869 224681 239897
rect 224709 239869 239979 239897
rect 240007 239869 240041 239897
rect 240069 239869 256437 239897
rect 256465 239869 256499 239897
rect 256527 239869 256561 239897
rect 256589 239869 256623 239897
rect 256651 239869 265437 239897
rect 265465 239869 265499 239897
rect 265527 239869 265561 239897
rect 265589 239869 265623 239897
rect 265651 239869 274437 239897
rect 274465 239869 274499 239897
rect 274527 239869 274561 239897
rect 274589 239869 274623 239897
rect 274651 239869 283437 239897
rect 283465 239869 283499 239897
rect 283527 239869 283561 239897
rect 283589 239869 283623 239897
rect 283651 239869 292437 239897
rect 292465 239869 292499 239897
rect 292527 239869 292561 239897
rect 292589 239869 292623 239897
rect 292651 239869 299736 239897
rect 299764 239869 299798 239897
rect 299826 239869 299860 239897
rect 299888 239869 299922 239897
rect 299950 239869 299998 239897
rect -6 239835 299998 239869
rect -6 239807 42 239835
rect 70 239807 104 239835
rect 132 239807 166 239835
rect 194 239807 228 239835
rect 256 239807 4437 239835
rect 4465 239807 4499 239835
rect 4527 239807 4561 239835
rect 4589 239807 4623 239835
rect 4651 239807 13437 239835
rect 13465 239807 13499 239835
rect 13527 239807 13561 239835
rect 13589 239807 13623 239835
rect 13651 239807 22437 239835
rect 22465 239807 22499 239835
rect 22527 239807 22561 239835
rect 22589 239807 22623 239835
rect 22651 239807 24939 239835
rect 24967 239807 25001 239835
rect 25029 239807 31437 239835
rect 31465 239807 31499 239835
rect 31527 239807 31561 239835
rect 31589 239807 31623 239835
rect 31651 239807 40299 239835
rect 40327 239807 40361 239835
rect 40389 239807 55659 239835
rect 55687 239807 55721 239835
rect 55749 239807 71019 239835
rect 71047 239807 71081 239835
rect 71109 239807 86379 239835
rect 86407 239807 86441 239835
rect 86469 239807 101739 239835
rect 101767 239807 101801 239835
rect 101829 239807 117099 239835
rect 117127 239807 117161 239835
rect 117189 239807 132459 239835
rect 132487 239807 132521 239835
rect 132549 239807 147819 239835
rect 147847 239807 147881 239835
rect 147909 239807 163179 239835
rect 163207 239807 163241 239835
rect 163269 239807 178539 239835
rect 178567 239807 178601 239835
rect 178629 239807 193899 239835
rect 193927 239807 193961 239835
rect 193989 239807 209259 239835
rect 209287 239807 209321 239835
rect 209349 239807 224619 239835
rect 224647 239807 224681 239835
rect 224709 239807 239979 239835
rect 240007 239807 240041 239835
rect 240069 239807 256437 239835
rect 256465 239807 256499 239835
rect 256527 239807 256561 239835
rect 256589 239807 256623 239835
rect 256651 239807 265437 239835
rect 265465 239807 265499 239835
rect 265527 239807 265561 239835
rect 265589 239807 265623 239835
rect 265651 239807 274437 239835
rect 274465 239807 274499 239835
rect 274527 239807 274561 239835
rect 274589 239807 274623 239835
rect 274651 239807 283437 239835
rect 283465 239807 283499 239835
rect 283527 239807 283561 239835
rect 283589 239807 283623 239835
rect 283651 239807 292437 239835
rect 292465 239807 292499 239835
rect 292527 239807 292561 239835
rect 292589 239807 292623 239835
rect 292651 239807 299736 239835
rect 299764 239807 299798 239835
rect 299826 239807 299860 239835
rect 299888 239807 299922 239835
rect 299950 239807 299998 239835
rect -6 239773 299998 239807
rect -6 239745 42 239773
rect 70 239745 104 239773
rect 132 239745 166 239773
rect 194 239745 228 239773
rect 256 239745 4437 239773
rect 4465 239745 4499 239773
rect 4527 239745 4561 239773
rect 4589 239745 4623 239773
rect 4651 239745 13437 239773
rect 13465 239745 13499 239773
rect 13527 239745 13561 239773
rect 13589 239745 13623 239773
rect 13651 239745 22437 239773
rect 22465 239745 22499 239773
rect 22527 239745 22561 239773
rect 22589 239745 22623 239773
rect 22651 239745 24939 239773
rect 24967 239745 25001 239773
rect 25029 239745 31437 239773
rect 31465 239745 31499 239773
rect 31527 239745 31561 239773
rect 31589 239745 31623 239773
rect 31651 239745 40299 239773
rect 40327 239745 40361 239773
rect 40389 239745 55659 239773
rect 55687 239745 55721 239773
rect 55749 239745 71019 239773
rect 71047 239745 71081 239773
rect 71109 239745 86379 239773
rect 86407 239745 86441 239773
rect 86469 239745 101739 239773
rect 101767 239745 101801 239773
rect 101829 239745 117099 239773
rect 117127 239745 117161 239773
rect 117189 239745 132459 239773
rect 132487 239745 132521 239773
rect 132549 239745 147819 239773
rect 147847 239745 147881 239773
rect 147909 239745 163179 239773
rect 163207 239745 163241 239773
rect 163269 239745 178539 239773
rect 178567 239745 178601 239773
rect 178629 239745 193899 239773
rect 193927 239745 193961 239773
rect 193989 239745 209259 239773
rect 209287 239745 209321 239773
rect 209349 239745 224619 239773
rect 224647 239745 224681 239773
rect 224709 239745 239979 239773
rect 240007 239745 240041 239773
rect 240069 239745 256437 239773
rect 256465 239745 256499 239773
rect 256527 239745 256561 239773
rect 256589 239745 256623 239773
rect 256651 239745 265437 239773
rect 265465 239745 265499 239773
rect 265527 239745 265561 239773
rect 265589 239745 265623 239773
rect 265651 239745 274437 239773
rect 274465 239745 274499 239773
rect 274527 239745 274561 239773
rect 274589 239745 274623 239773
rect 274651 239745 283437 239773
rect 283465 239745 283499 239773
rect 283527 239745 283561 239773
rect 283589 239745 283623 239773
rect 283651 239745 292437 239773
rect 292465 239745 292499 239773
rect 292527 239745 292561 239773
rect 292589 239745 292623 239773
rect 292651 239745 299736 239773
rect 299764 239745 299798 239773
rect 299826 239745 299860 239773
rect 299888 239745 299922 239773
rect 299950 239745 299998 239773
rect -6 239697 299998 239745
rect -6 236959 299998 237007
rect -6 236931 522 236959
rect 550 236931 584 236959
rect 612 236931 646 236959
rect 674 236931 708 236959
rect 736 236931 2577 236959
rect 2605 236931 2639 236959
rect 2667 236931 2701 236959
rect 2729 236931 2763 236959
rect 2791 236931 11577 236959
rect 11605 236931 11639 236959
rect 11667 236931 11701 236959
rect 11729 236931 11763 236959
rect 11791 236931 17259 236959
rect 17287 236931 17321 236959
rect 17349 236931 20577 236959
rect 20605 236931 20639 236959
rect 20667 236931 20701 236959
rect 20729 236931 20763 236959
rect 20791 236931 29577 236959
rect 29605 236931 29639 236959
rect 29667 236931 29701 236959
rect 29729 236931 29763 236959
rect 29791 236931 32619 236959
rect 32647 236931 32681 236959
rect 32709 236931 47979 236959
rect 48007 236931 48041 236959
rect 48069 236931 63339 236959
rect 63367 236931 63401 236959
rect 63429 236931 78699 236959
rect 78727 236931 78761 236959
rect 78789 236931 94059 236959
rect 94087 236931 94121 236959
rect 94149 236931 109419 236959
rect 109447 236931 109481 236959
rect 109509 236931 124779 236959
rect 124807 236931 124841 236959
rect 124869 236931 140139 236959
rect 140167 236931 140201 236959
rect 140229 236931 155499 236959
rect 155527 236931 155561 236959
rect 155589 236931 170859 236959
rect 170887 236931 170921 236959
rect 170949 236931 186219 236959
rect 186247 236931 186281 236959
rect 186309 236931 201579 236959
rect 201607 236931 201641 236959
rect 201669 236931 216939 236959
rect 216967 236931 217001 236959
rect 217029 236931 232299 236959
rect 232327 236931 232361 236959
rect 232389 236931 247659 236959
rect 247687 236931 247721 236959
rect 247749 236931 254577 236959
rect 254605 236931 254639 236959
rect 254667 236931 254701 236959
rect 254729 236931 254763 236959
rect 254791 236931 263577 236959
rect 263605 236931 263639 236959
rect 263667 236931 263701 236959
rect 263729 236931 263763 236959
rect 263791 236931 272577 236959
rect 272605 236931 272639 236959
rect 272667 236931 272701 236959
rect 272729 236931 272763 236959
rect 272791 236931 281577 236959
rect 281605 236931 281639 236959
rect 281667 236931 281701 236959
rect 281729 236931 281763 236959
rect 281791 236931 290577 236959
rect 290605 236931 290639 236959
rect 290667 236931 290701 236959
rect 290729 236931 290763 236959
rect 290791 236931 299256 236959
rect 299284 236931 299318 236959
rect 299346 236931 299380 236959
rect 299408 236931 299442 236959
rect 299470 236931 299998 236959
rect -6 236897 299998 236931
rect -6 236869 522 236897
rect 550 236869 584 236897
rect 612 236869 646 236897
rect 674 236869 708 236897
rect 736 236869 2577 236897
rect 2605 236869 2639 236897
rect 2667 236869 2701 236897
rect 2729 236869 2763 236897
rect 2791 236869 11577 236897
rect 11605 236869 11639 236897
rect 11667 236869 11701 236897
rect 11729 236869 11763 236897
rect 11791 236869 17259 236897
rect 17287 236869 17321 236897
rect 17349 236869 20577 236897
rect 20605 236869 20639 236897
rect 20667 236869 20701 236897
rect 20729 236869 20763 236897
rect 20791 236869 29577 236897
rect 29605 236869 29639 236897
rect 29667 236869 29701 236897
rect 29729 236869 29763 236897
rect 29791 236869 32619 236897
rect 32647 236869 32681 236897
rect 32709 236869 47979 236897
rect 48007 236869 48041 236897
rect 48069 236869 63339 236897
rect 63367 236869 63401 236897
rect 63429 236869 78699 236897
rect 78727 236869 78761 236897
rect 78789 236869 94059 236897
rect 94087 236869 94121 236897
rect 94149 236869 109419 236897
rect 109447 236869 109481 236897
rect 109509 236869 124779 236897
rect 124807 236869 124841 236897
rect 124869 236869 140139 236897
rect 140167 236869 140201 236897
rect 140229 236869 155499 236897
rect 155527 236869 155561 236897
rect 155589 236869 170859 236897
rect 170887 236869 170921 236897
rect 170949 236869 186219 236897
rect 186247 236869 186281 236897
rect 186309 236869 201579 236897
rect 201607 236869 201641 236897
rect 201669 236869 216939 236897
rect 216967 236869 217001 236897
rect 217029 236869 232299 236897
rect 232327 236869 232361 236897
rect 232389 236869 247659 236897
rect 247687 236869 247721 236897
rect 247749 236869 254577 236897
rect 254605 236869 254639 236897
rect 254667 236869 254701 236897
rect 254729 236869 254763 236897
rect 254791 236869 263577 236897
rect 263605 236869 263639 236897
rect 263667 236869 263701 236897
rect 263729 236869 263763 236897
rect 263791 236869 272577 236897
rect 272605 236869 272639 236897
rect 272667 236869 272701 236897
rect 272729 236869 272763 236897
rect 272791 236869 281577 236897
rect 281605 236869 281639 236897
rect 281667 236869 281701 236897
rect 281729 236869 281763 236897
rect 281791 236869 290577 236897
rect 290605 236869 290639 236897
rect 290667 236869 290701 236897
rect 290729 236869 290763 236897
rect 290791 236869 299256 236897
rect 299284 236869 299318 236897
rect 299346 236869 299380 236897
rect 299408 236869 299442 236897
rect 299470 236869 299998 236897
rect -6 236835 299998 236869
rect -6 236807 522 236835
rect 550 236807 584 236835
rect 612 236807 646 236835
rect 674 236807 708 236835
rect 736 236807 2577 236835
rect 2605 236807 2639 236835
rect 2667 236807 2701 236835
rect 2729 236807 2763 236835
rect 2791 236807 11577 236835
rect 11605 236807 11639 236835
rect 11667 236807 11701 236835
rect 11729 236807 11763 236835
rect 11791 236807 17259 236835
rect 17287 236807 17321 236835
rect 17349 236807 20577 236835
rect 20605 236807 20639 236835
rect 20667 236807 20701 236835
rect 20729 236807 20763 236835
rect 20791 236807 29577 236835
rect 29605 236807 29639 236835
rect 29667 236807 29701 236835
rect 29729 236807 29763 236835
rect 29791 236807 32619 236835
rect 32647 236807 32681 236835
rect 32709 236807 47979 236835
rect 48007 236807 48041 236835
rect 48069 236807 63339 236835
rect 63367 236807 63401 236835
rect 63429 236807 78699 236835
rect 78727 236807 78761 236835
rect 78789 236807 94059 236835
rect 94087 236807 94121 236835
rect 94149 236807 109419 236835
rect 109447 236807 109481 236835
rect 109509 236807 124779 236835
rect 124807 236807 124841 236835
rect 124869 236807 140139 236835
rect 140167 236807 140201 236835
rect 140229 236807 155499 236835
rect 155527 236807 155561 236835
rect 155589 236807 170859 236835
rect 170887 236807 170921 236835
rect 170949 236807 186219 236835
rect 186247 236807 186281 236835
rect 186309 236807 201579 236835
rect 201607 236807 201641 236835
rect 201669 236807 216939 236835
rect 216967 236807 217001 236835
rect 217029 236807 232299 236835
rect 232327 236807 232361 236835
rect 232389 236807 247659 236835
rect 247687 236807 247721 236835
rect 247749 236807 254577 236835
rect 254605 236807 254639 236835
rect 254667 236807 254701 236835
rect 254729 236807 254763 236835
rect 254791 236807 263577 236835
rect 263605 236807 263639 236835
rect 263667 236807 263701 236835
rect 263729 236807 263763 236835
rect 263791 236807 272577 236835
rect 272605 236807 272639 236835
rect 272667 236807 272701 236835
rect 272729 236807 272763 236835
rect 272791 236807 281577 236835
rect 281605 236807 281639 236835
rect 281667 236807 281701 236835
rect 281729 236807 281763 236835
rect 281791 236807 290577 236835
rect 290605 236807 290639 236835
rect 290667 236807 290701 236835
rect 290729 236807 290763 236835
rect 290791 236807 299256 236835
rect 299284 236807 299318 236835
rect 299346 236807 299380 236835
rect 299408 236807 299442 236835
rect 299470 236807 299998 236835
rect -6 236773 299998 236807
rect -6 236745 522 236773
rect 550 236745 584 236773
rect 612 236745 646 236773
rect 674 236745 708 236773
rect 736 236745 2577 236773
rect 2605 236745 2639 236773
rect 2667 236745 2701 236773
rect 2729 236745 2763 236773
rect 2791 236745 11577 236773
rect 11605 236745 11639 236773
rect 11667 236745 11701 236773
rect 11729 236745 11763 236773
rect 11791 236745 17259 236773
rect 17287 236745 17321 236773
rect 17349 236745 20577 236773
rect 20605 236745 20639 236773
rect 20667 236745 20701 236773
rect 20729 236745 20763 236773
rect 20791 236745 29577 236773
rect 29605 236745 29639 236773
rect 29667 236745 29701 236773
rect 29729 236745 29763 236773
rect 29791 236745 32619 236773
rect 32647 236745 32681 236773
rect 32709 236745 47979 236773
rect 48007 236745 48041 236773
rect 48069 236745 63339 236773
rect 63367 236745 63401 236773
rect 63429 236745 78699 236773
rect 78727 236745 78761 236773
rect 78789 236745 94059 236773
rect 94087 236745 94121 236773
rect 94149 236745 109419 236773
rect 109447 236745 109481 236773
rect 109509 236745 124779 236773
rect 124807 236745 124841 236773
rect 124869 236745 140139 236773
rect 140167 236745 140201 236773
rect 140229 236745 155499 236773
rect 155527 236745 155561 236773
rect 155589 236745 170859 236773
rect 170887 236745 170921 236773
rect 170949 236745 186219 236773
rect 186247 236745 186281 236773
rect 186309 236745 201579 236773
rect 201607 236745 201641 236773
rect 201669 236745 216939 236773
rect 216967 236745 217001 236773
rect 217029 236745 232299 236773
rect 232327 236745 232361 236773
rect 232389 236745 247659 236773
rect 247687 236745 247721 236773
rect 247749 236745 254577 236773
rect 254605 236745 254639 236773
rect 254667 236745 254701 236773
rect 254729 236745 254763 236773
rect 254791 236745 263577 236773
rect 263605 236745 263639 236773
rect 263667 236745 263701 236773
rect 263729 236745 263763 236773
rect 263791 236745 272577 236773
rect 272605 236745 272639 236773
rect 272667 236745 272701 236773
rect 272729 236745 272763 236773
rect 272791 236745 281577 236773
rect 281605 236745 281639 236773
rect 281667 236745 281701 236773
rect 281729 236745 281763 236773
rect 281791 236745 290577 236773
rect 290605 236745 290639 236773
rect 290667 236745 290701 236773
rect 290729 236745 290763 236773
rect 290791 236745 299256 236773
rect 299284 236745 299318 236773
rect 299346 236745 299380 236773
rect 299408 236745 299442 236773
rect 299470 236745 299998 236773
rect -6 236697 299998 236745
rect -6 230959 299998 231007
rect -6 230931 42 230959
rect 70 230931 104 230959
rect 132 230931 166 230959
rect 194 230931 228 230959
rect 256 230931 4437 230959
rect 4465 230931 4499 230959
rect 4527 230931 4561 230959
rect 4589 230931 4623 230959
rect 4651 230931 13437 230959
rect 13465 230931 13499 230959
rect 13527 230931 13561 230959
rect 13589 230931 13623 230959
rect 13651 230931 22437 230959
rect 22465 230931 22499 230959
rect 22527 230931 22561 230959
rect 22589 230931 22623 230959
rect 22651 230931 24939 230959
rect 24967 230931 25001 230959
rect 25029 230931 31437 230959
rect 31465 230931 31499 230959
rect 31527 230931 31561 230959
rect 31589 230931 31623 230959
rect 31651 230931 40299 230959
rect 40327 230931 40361 230959
rect 40389 230931 55659 230959
rect 55687 230931 55721 230959
rect 55749 230931 71019 230959
rect 71047 230931 71081 230959
rect 71109 230931 86379 230959
rect 86407 230931 86441 230959
rect 86469 230931 101739 230959
rect 101767 230931 101801 230959
rect 101829 230931 117099 230959
rect 117127 230931 117161 230959
rect 117189 230931 132459 230959
rect 132487 230931 132521 230959
rect 132549 230931 147819 230959
rect 147847 230931 147881 230959
rect 147909 230931 163179 230959
rect 163207 230931 163241 230959
rect 163269 230931 178539 230959
rect 178567 230931 178601 230959
rect 178629 230931 193899 230959
rect 193927 230931 193961 230959
rect 193989 230931 209259 230959
rect 209287 230931 209321 230959
rect 209349 230931 224619 230959
rect 224647 230931 224681 230959
rect 224709 230931 239979 230959
rect 240007 230931 240041 230959
rect 240069 230931 256437 230959
rect 256465 230931 256499 230959
rect 256527 230931 256561 230959
rect 256589 230931 256623 230959
rect 256651 230931 265437 230959
rect 265465 230931 265499 230959
rect 265527 230931 265561 230959
rect 265589 230931 265623 230959
rect 265651 230931 274437 230959
rect 274465 230931 274499 230959
rect 274527 230931 274561 230959
rect 274589 230931 274623 230959
rect 274651 230931 283437 230959
rect 283465 230931 283499 230959
rect 283527 230931 283561 230959
rect 283589 230931 283623 230959
rect 283651 230931 292437 230959
rect 292465 230931 292499 230959
rect 292527 230931 292561 230959
rect 292589 230931 292623 230959
rect 292651 230931 299736 230959
rect 299764 230931 299798 230959
rect 299826 230931 299860 230959
rect 299888 230931 299922 230959
rect 299950 230931 299998 230959
rect -6 230897 299998 230931
rect -6 230869 42 230897
rect 70 230869 104 230897
rect 132 230869 166 230897
rect 194 230869 228 230897
rect 256 230869 4437 230897
rect 4465 230869 4499 230897
rect 4527 230869 4561 230897
rect 4589 230869 4623 230897
rect 4651 230869 13437 230897
rect 13465 230869 13499 230897
rect 13527 230869 13561 230897
rect 13589 230869 13623 230897
rect 13651 230869 22437 230897
rect 22465 230869 22499 230897
rect 22527 230869 22561 230897
rect 22589 230869 22623 230897
rect 22651 230869 24939 230897
rect 24967 230869 25001 230897
rect 25029 230869 31437 230897
rect 31465 230869 31499 230897
rect 31527 230869 31561 230897
rect 31589 230869 31623 230897
rect 31651 230869 40299 230897
rect 40327 230869 40361 230897
rect 40389 230869 55659 230897
rect 55687 230869 55721 230897
rect 55749 230869 71019 230897
rect 71047 230869 71081 230897
rect 71109 230869 86379 230897
rect 86407 230869 86441 230897
rect 86469 230869 101739 230897
rect 101767 230869 101801 230897
rect 101829 230869 117099 230897
rect 117127 230869 117161 230897
rect 117189 230869 132459 230897
rect 132487 230869 132521 230897
rect 132549 230869 147819 230897
rect 147847 230869 147881 230897
rect 147909 230869 163179 230897
rect 163207 230869 163241 230897
rect 163269 230869 178539 230897
rect 178567 230869 178601 230897
rect 178629 230869 193899 230897
rect 193927 230869 193961 230897
rect 193989 230869 209259 230897
rect 209287 230869 209321 230897
rect 209349 230869 224619 230897
rect 224647 230869 224681 230897
rect 224709 230869 239979 230897
rect 240007 230869 240041 230897
rect 240069 230869 256437 230897
rect 256465 230869 256499 230897
rect 256527 230869 256561 230897
rect 256589 230869 256623 230897
rect 256651 230869 265437 230897
rect 265465 230869 265499 230897
rect 265527 230869 265561 230897
rect 265589 230869 265623 230897
rect 265651 230869 274437 230897
rect 274465 230869 274499 230897
rect 274527 230869 274561 230897
rect 274589 230869 274623 230897
rect 274651 230869 283437 230897
rect 283465 230869 283499 230897
rect 283527 230869 283561 230897
rect 283589 230869 283623 230897
rect 283651 230869 292437 230897
rect 292465 230869 292499 230897
rect 292527 230869 292561 230897
rect 292589 230869 292623 230897
rect 292651 230869 299736 230897
rect 299764 230869 299798 230897
rect 299826 230869 299860 230897
rect 299888 230869 299922 230897
rect 299950 230869 299998 230897
rect -6 230835 299998 230869
rect -6 230807 42 230835
rect 70 230807 104 230835
rect 132 230807 166 230835
rect 194 230807 228 230835
rect 256 230807 4437 230835
rect 4465 230807 4499 230835
rect 4527 230807 4561 230835
rect 4589 230807 4623 230835
rect 4651 230807 13437 230835
rect 13465 230807 13499 230835
rect 13527 230807 13561 230835
rect 13589 230807 13623 230835
rect 13651 230807 22437 230835
rect 22465 230807 22499 230835
rect 22527 230807 22561 230835
rect 22589 230807 22623 230835
rect 22651 230807 24939 230835
rect 24967 230807 25001 230835
rect 25029 230807 31437 230835
rect 31465 230807 31499 230835
rect 31527 230807 31561 230835
rect 31589 230807 31623 230835
rect 31651 230807 40299 230835
rect 40327 230807 40361 230835
rect 40389 230807 55659 230835
rect 55687 230807 55721 230835
rect 55749 230807 71019 230835
rect 71047 230807 71081 230835
rect 71109 230807 86379 230835
rect 86407 230807 86441 230835
rect 86469 230807 101739 230835
rect 101767 230807 101801 230835
rect 101829 230807 117099 230835
rect 117127 230807 117161 230835
rect 117189 230807 132459 230835
rect 132487 230807 132521 230835
rect 132549 230807 147819 230835
rect 147847 230807 147881 230835
rect 147909 230807 163179 230835
rect 163207 230807 163241 230835
rect 163269 230807 178539 230835
rect 178567 230807 178601 230835
rect 178629 230807 193899 230835
rect 193927 230807 193961 230835
rect 193989 230807 209259 230835
rect 209287 230807 209321 230835
rect 209349 230807 224619 230835
rect 224647 230807 224681 230835
rect 224709 230807 239979 230835
rect 240007 230807 240041 230835
rect 240069 230807 256437 230835
rect 256465 230807 256499 230835
rect 256527 230807 256561 230835
rect 256589 230807 256623 230835
rect 256651 230807 265437 230835
rect 265465 230807 265499 230835
rect 265527 230807 265561 230835
rect 265589 230807 265623 230835
rect 265651 230807 274437 230835
rect 274465 230807 274499 230835
rect 274527 230807 274561 230835
rect 274589 230807 274623 230835
rect 274651 230807 283437 230835
rect 283465 230807 283499 230835
rect 283527 230807 283561 230835
rect 283589 230807 283623 230835
rect 283651 230807 292437 230835
rect 292465 230807 292499 230835
rect 292527 230807 292561 230835
rect 292589 230807 292623 230835
rect 292651 230807 299736 230835
rect 299764 230807 299798 230835
rect 299826 230807 299860 230835
rect 299888 230807 299922 230835
rect 299950 230807 299998 230835
rect -6 230773 299998 230807
rect -6 230745 42 230773
rect 70 230745 104 230773
rect 132 230745 166 230773
rect 194 230745 228 230773
rect 256 230745 4437 230773
rect 4465 230745 4499 230773
rect 4527 230745 4561 230773
rect 4589 230745 4623 230773
rect 4651 230745 13437 230773
rect 13465 230745 13499 230773
rect 13527 230745 13561 230773
rect 13589 230745 13623 230773
rect 13651 230745 22437 230773
rect 22465 230745 22499 230773
rect 22527 230745 22561 230773
rect 22589 230745 22623 230773
rect 22651 230745 24939 230773
rect 24967 230745 25001 230773
rect 25029 230745 31437 230773
rect 31465 230745 31499 230773
rect 31527 230745 31561 230773
rect 31589 230745 31623 230773
rect 31651 230745 40299 230773
rect 40327 230745 40361 230773
rect 40389 230745 55659 230773
rect 55687 230745 55721 230773
rect 55749 230745 71019 230773
rect 71047 230745 71081 230773
rect 71109 230745 86379 230773
rect 86407 230745 86441 230773
rect 86469 230745 101739 230773
rect 101767 230745 101801 230773
rect 101829 230745 117099 230773
rect 117127 230745 117161 230773
rect 117189 230745 132459 230773
rect 132487 230745 132521 230773
rect 132549 230745 147819 230773
rect 147847 230745 147881 230773
rect 147909 230745 163179 230773
rect 163207 230745 163241 230773
rect 163269 230745 178539 230773
rect 178567 230745 178601 230773
rect 178629 230745 193899 230773
rect 193927 230745 193961 230773
rect 193989 230745 209259 230773
rect 209287 230745 209321 230773
rect 209349 230745 224619 230773
rect 224647 230745 224681 230773
rect 224709 230745 239979 230773
rect 240007 230745 240041 230773
rect 240069 230745 256437 230773
rect 256465 230745 256499 230773
rect 256527 230745 256561 230773
rect 256589 230745 256623 230773
rect 256651 230745 265437 230773
rect 265465 230745 265499 230773
rect 265527 230745 265561 230773
rect 265589 230745 265623 230773
rect 265651 230745 274437 230773
rect 274465 230745 274499 230773
rect 274527 230745 274561 230773
rect 274589 230745 274623 230773
rect 274651 230745 283437 230773
rect 283465 230745 283499 230773
rect 283527 230745 283561 230773
rect 283589 230745 283623 230773
rect 283651 230745 292437 230773
rect 292465 230745 292499 230773
rect 292527 230745 292561 230773
rect 292589 230745 292623 230773
rect 292651 230745 299736 230773
rect 299764 230745 299798 230773
rect 299826 230745 299860 230773
rect 299888 230745 299922 230773
rect 299950 230745 299998 230773
rect -6 230697 299998 230745
rect -6 227959 299998 228007
rect -6 227931 522 227959
rect 550 227931 584 227959
rect 612 227931 646 227959
rect 674 227931 708 227959
rect 736 227931 2577 227959
rect 2605 227931 2639 227959
rect 2667 227931 2701 227959
rect 2729 227931 2763 227959
rect 2791 227931 11577 227959
rect 11605 227931 11639 227959
rect 11667 227931 11701 227959
rect 11729 227931 11763 227959
rect 11791 227931 17259 227959
rect 17287 227931 17321 227959
rect 17349 227931 20577 227959
rect 20605 227931 20639 227959
rect 20667 227931 20701 227959
rect 20729 227931 20763 227959
rect 20791 227931 29577 227959
rect 29605 227931 29639 227959
rect 29667 227931 29701 227959
rect 29729 227931 29763 227959
rect 29791 227931 32619 227959
rect 32647 227931 32681 227959
rect 32709 227931 47979 227959
rect 48007 227931 48041 227959
rect 48069 227931 63339 227959
rect 63367 227931 63401 227959
rect 63429 227931 78699 227959
rect 78727 227931 78761 227959
rect 78789 227931 94059 227959
rect 94087 227931 94121 227959
rect 94149 227931 109419 227959
rect 109447 227931 109481 227959
rect 109509 227931 124779 227959
rect 124807 227931 124841 227959
rect 124869 227931 140139 227959
rect 140167 227931 140201 227959
rect 140229 227931 155499 227959
rect 155527 227931 155561 227959
rect 155589 227931 170859 227959
rect 170887 227931 170921 227959
rect 170949 227931 186219 227959
rect 186247 227931 186281 227959
rect 186309 227931 201579 227959
rect 201607 227931 201641 227959
rect 201669 227931 216939 227959
rect 216967 227931 217001 227959
rect 217029 227931 232299 227959
rect 232327 227931 232361 227959
rect 232389 227931 247659 227959
rect 247687 227931 247721 227959
rect 247749 227931 254577 227959
rect 254605 227931 254639 227959
rect 254667 227931 254701 227959
rect 254729 227931 254763 227959
rect 254791 227931 263577 227959
rect 263605 227931 263639 227959
rect 263667 227931 263701 227959
rect 263729 227931 263763 227959
rect 263791 227931 272577 227959
rect 272605 227931 272639 227959
rect 272667 227931 272701 227959
rect 272729 227931 272763 227959
rect 272791 227931 281577 227959
rect 281605 227931 281639 227959
rect 281667 227931 281701 227959
rect 281729 227931 281763 227959
rect 281791 227931 290577 227959
rect 290605 227931 290639 227959
rect 290667 227931 290701 227959
rect 290729 227931 290763 227959
rect 290791 227931 299256 227959
rect 299284 227931 299318 227959
rect 299346 227931 299380 227959
rect 299408 227931 299442 227959
rect 299470 227931 299998 227959
rect -6 227897 299998 227931
rect -6 227869 522 227897
rect 550 227869 584 227897
rect 612 227869 646 227897
rect 674 227869 708 227897
rect 736 227869 2577 227897
rect 2605 227869 2639 227897
rect 2667 227869 2701 227897
rect 2729 227869 2763 227897
rect 2791 227869 11577 227897
rect 11605 227869 11639 227897
rect 11667 227869 11701 227897
rect 11729 227869 11763 227897
rect 11791 227869 17259 227897
rect 17287 227869 17321 227897
rect 17349 227869 20577 227897
rect 20605 227869 20639 227897
rect 20667 227869 20701 227897
rect 20729 227869 20763 227897
rect 20791 227869 29577 227897
rect 29605 227869 29639 227897
rect 29667 227869 29701 227897
rect 29729 227869 29763 227897
rect 29791 227869 32619 227897
rect 32647 227869 32681 227897
rect 32709 227869 47979 227897
rect 48007 227869 48041 227897
rect 48069 227869 63339 227897
rect 63367 227869 63401 227897
rect 63429 227869 78699 227897
rect 78727 227869 78761 227897
rect 78789 227869 94059 227897
rect 94087 227869 94121 227897
rect 94149 227869 109419 227897
rect 109447 227869 109481 227897
rect 109509 227869 124779 227897
rect 124807 227869 124841 227897
rect 124869 227869 140139 227897
rect 140167 227869 140201 227897
rect 140229 227869 155499 227897
rect 155527 227869 155561 227897
rect 155589 227869 170859 227897
rect 170887 227869 170921 227897
rect 170949 227869 186219 227897
rect 186247 227869 186281 227897
rect 186309 227869 201579 227897
rect 201607 227869 201641 227897
rect 201669 227869 216939 227897
rect 216967 227869 217001 227897
rect 217029 227869 232299 227897
rect 232327 227869 232361 227897
rect 232389 227869 247659 227897
rect 247687 227869 247721 227897
rect 247749 227869 254577 227897
rect 254605 227869 254639 227897
rect 254667 227869 254701 227897
rect 254729 227869 254763 227897
rect 254791 227869 263577 227897
rect 263605 227869 263639 227897
rect 263667 227869 263701 227897
rect 263729 227869 263763 227897
rect 263791 227869 272577 227897
rect 272605 227869 272639 227897
rect 272667 227869 272701 227897
rect 272729 227869 272763 227897
rect 272791 227869 281577 227897
rect 281605 227869 281639 227897
rect 281667 227869 281701 227897
rect 281729 227869 281763 227897
rect 281791 227869 290577 227897
rect 290605 227869 290639 227897
rect 290667 227869 290701 227897
rect 290729 227869 290763 227897
rect 290791 227869 299256 227897
rect 299284 227869 299318 227897
rect 299346 227869 299380 227897
rect 299408 227869 299442 227897
rect 299470 227869 299998 227897
rect -6 227835 299998 227869
rect -6 227807 522 227835
rect 550 227807 584 227835
rect 612 227807 646 227835
rect 674 227807 708 227835
rect 736 227807 2577 227835
rect 2605 227807 2639 227835
rect 2667 227807 2701 227835
rect 2729 227807 2763 227835
rect 2791 227807 11577 227835
rect 11605 227807 11639 227835
rect 11667 227807 11701 227835
rect 11729 227807 11763 227835
rect 11791 227807 17259 227835
rect 17287 227807 17321 227835
rect 17349 227807 20577 227835
rect 20605 227807 20639 227835
rect 20667 227807 20701 227835
rect 20729 227807 20763 227835
rect 20791 227807 29577 227835
rect 29605 227807 29639 227835
rect 29667 227807 29701 227835
rect 29729 227807 29763 227835
rect 29791 227807 32619 227835
rect 32647 227807 32681 227835
rect 32709 227807 47979 227835
rect 48007 227807 48041 227835
rect 48069 227807 63339 227835
rect 63367 227807 63401 227835
rect 63429 227807 78699 227835
rect 78727 227807 78761 227835
rect 78789 227807 94059 227835
rect 94087 227807 94121 227835
rect 94149 227807 109419 227835
rect 109447 227807 109481 227835
rect 109509 227807 124779 227835
rect 124807 227807 124841 227835
rect 124869 227807 140139 227835
rect 140167 227807 140201 227835
rect 140229 227807 155499 227835
rect 155527 227807 155561 227835
rect 155589 227807 170859 227835
rect 170887 227807 170921 227835
rect 170949 227807 186219 227835
rect 186247 227807 186281 227835
rect 186309 227807 201579 227835
rect 201607 227807 201641 227835
rect 201669 227807 216939 227835
rect 216967 227807 217001 227835
rect 217029 227807 232299 227835
rect 232327 227807 232361 227835
rect 232389 227807 247659 227835
rect 247687 227807 247721 227835
rect 247749 227807 254577 227835
rect 254605 227807 254639 227835
rect 254667 227807 254701 227835
rect 254729 227807 254763 227835
rect 254791 227807 263577 227835
rect 263605 227807 263639 227835
rect 263667 227807 263701 227835
rect 263729 227807 263763 227835
rect 263791 227807 272577 227835
rect 272605 227807 272639 227835
rect 272667 227807 272701 227835
rect 272729 227807 272763 227835
rect 272791 227807 281577 227835
rect 281605 227807 281639 227835
rect 281667 227807 281701 227835
rect 281729 227807 281763 227835
rect 281791 227807 290577 227835
rect 290605 227807 290639 227835
rect 290667 227807 290701 227835
rect 290729 227807 290763 227835
rect 290791 227807 299256 227835
rect 299284 227807 299318 227835
rect 299346 227807 299380 227835
rect 299408 227807 299442 227835
rect 299470 227807 299998 227835
rect -6 227773 299998 227807
rect -6 227745 522 227773
rect 550 227745 584 227773
rect 612 227745 646 227773
rect 674 227745 708 227773
rect 736 227745 2577 227773
rect 2605 227745 2639 227773
rect 2667 227745 2701 227773
rect 2729 227745 2763 227773
rect 2791 227745 11577 227773
rect 11605 227745 11639 227773
rect 11667 227745 11701 227773
rect 11729 227745 11763 227773
rect 11791 227745 17259 227773
rect 17287 227745 17321 227773
rect 17349 227745 20577 227773
rect 20605 227745 20639 227773
rect 20667 227745 20701 227773
rect 20729 227745 20763 227773
rect 20791 227745 29577 227773
rect 29605 227745 29639 227773
rect 29667 227745 29701 227773
rect 29729 227745 29763 227773
rect 29791 227745 32619 227773
rect 32647 227745 32681 227773
rect 32709 227745 47979 227773
rect 48007 227745 48041 227773
rect 48069 227745 63339 227773
rect 63367 227745 63401 227773
rect 63429 227745 78699 227773
rect 78727 227745 78761 227773
rect 78789 227745 94059 227773
rect 94087 227745 94121 227773
rect 94149 227745 109419 227773
rect 109447 227745 109481 227773
rect 109509 227745 124779 227773
rect 124807 227745 124841 227773
rect 124869 227745 140139 227773
rect 140167 227745 140201 227773
rect 140229 227745 155499 227773
rect 155527 227745 155561 227773
rect 155589 227745 170859 227773
rect 170887 227745 170921 227773
rect 170949 227745 186219 227773
rect 186247 227745 186281 227773
rect 186309 227745 201579 227773
rect 201607 227745 201641 227773
rect 201669 227745 216939 227773
rect 216967 227745 217001 227773
rect 217029 227745 232299 227773
rect 232327 227745 232361 227773
rect 232389 227745 247659 227773
rect 247687 227745 247721 227773
rect 247749 227745 254577 227773
rect 254605 227745 254639 227773
rect 254667 227745 254701 227773
rect 254729 227745 254763 227773
rect 254791 227745 263577 227773
rect 263605 227745 263639 227773
rect 263667 227745 263701 227773
rect 263729 227745 263763 227773
rect 263791 227745 272577 227773
rect 272605 227745 272639 227773
rect 272667 227745 272701 227773
rect 272729 227745 272763 227773
rect 272791 227745 281577 227773
rect 281605 227745 281639 227773
rect 281667 227745 281701 227773
rect 281729 227745 281763 227773
rect 281791 227745 290577 227773
rect 290605 227745 290639 227773
rect 290667 227745 290701 227773
rect 290729 227745 290763 227773
rect 290791 227745 299256 227773
rect 299284 227745 299318 227773
rect 299346 227745 299380 227773
rect 299408 227745 299442 227773
rect 299470 227745 299998 227773
rect -6 227697 299998 227745
rect -6 221959 299998 222007
rect -6 221931 42 221959
rect 70 221931 104 221959
rect 132 221931 166 221959
rect 194 221931 228 221959
rect 256 221931 4437 221959
rect 4465 221931 4499 221959
rect 4527 221931 4561 221959
rect 4589 221931 4623 221959
rect 4651 221931 13437 221959
rect 13465 221931 13499 221959
rect 13527 221931 13561 221959
rect 13589 221931 13623 221959
rect 13651 221931 22437 221959
rect 22465 221931 22499 221959
rect 22527 221931 22561 221959
rect 22589 221931 22623 221959
rect 22651 221931 24939 221959
rect 24967 221931 25001 221959
rect 25029 221931 31437 221959
rect 31465 221931 31499 221959
rect 31527 221931 31561 221959
rect 31589 221931 31623 221959
rect 31651 221931 40299 221959
rect 40327 221931 40361 221959
rect 40389 221931 55659 221959
rect 55687 221931 55721 221959
rect 55749 221931 71019 221959
rect 71047 221931 71081 221959
rect 71109 221931 86379 221959
rect 86407 221931 86441 221959
rect 86469 221931 101739 221959
rect 101767 221931 101801 221959
rect 101829 221931 117099 221959
rect 117127 221931 117161 221959
rect 117189 221931 132459 221959
rect 132487 221931 132521 221959
rect 132549 221931 147819 221959
rect 147847 221931 147881 221959
rect 147909 221931 163179 221959
rect 163207 221931 163241 221959
rect 163269 221931 178539 221959
rect 178567 221931 178601 221959
rect 178629 221931 193899 221959
rect 193927 221931 193961 221959
rect 193989 221931 209259 221959
rect 209287 221931 209321 221959
rect 209349 221931 224619 221959
rect 224647 221931 224681 221959
rect 224709 221931 239979 221959
rect 240007 221931 240041 221959
rect 240069 221931 256437 221959
rect 256465 221931 256499 221959
rect 256527 221931 256561 221959
rect 256589 221931 256623 221959
rect 256651 221931 265437 221959
rect 265465 221931 265499 221959
rect 265527 221931 265561 221959
rect 265589 221931 265623 221959
rect 265651 221931 274437 221959
rect 274465 221931 274499 221959
rect 274527 221931 274561 221959
rect 274589 221931 274623 221959
rect 274651 221931 283437 221959
rect 283465 221931 283499 221959
rect 283527 221931 283561 221959
rect 283589 221931 283623 221959
rect 283651 221931 292437 221959
rect 292465 221931 292499 221959
rect 292527 221931 292561 221959
rect 292589 221931 292623 221959
rect 292651 221931 299736 221959
rect 299764 221931 299798 221959
rect 299826 221931 299860 221959
rect 299888 221931 299922 221959
rect 299950 221931 299998 221959
rect -6 221897 299998 221931
rect -6 221869 42 221897
rect 70 221869 104 221897
rect 132 221869 166 221897
rect 194 221869 228 221897
rect 256 221869 4437 221897
rect 4465 221869 4499 221897
rect 4527 221869 4561 221897
rect 4589 221869 4623 221897
rect 4651 221869 13437 221897
rect 13465 221869 13499 221897
rect 13527 221869 13561 221897
rect 13589 221869 13623 221897
rect 13651 221869 22437 221897
rect 22465 221869 22499 221897
rect 22527 221869 22561 221897
rect 22589 221869 22623 221897
rect 22651 221869 24939 221897
rect 24967 221869 25001 221897
rect 25029 221869 31437 221897
rect 31465 221869 31499 221897
rect 31527 221869 31561 221897
rect 31589 221869 31623 221897
rect 31651 221869 40299 221897
rect 40327 221869 40361 221897
rect 40389 221869 55659 221897
rect 55687 221869 55721 221897
rect 55749 221869 71019 221897
rect 71047 221869 71081 221897
rect 71109 221869 86379 221897
rect 86407 221869 86441 221897
rect 86469 221869 101739 221897
rect 101767 221869 101801 221897
rect 101829 221869 117099 221897
rect 117127 221869 117161 221897
rect 117189 221869 132459 221897
rect 132487 221869 132521 221897
rect 132549 221869 147819 221897
rect 147847 221869 147881 221897
rect 147909 221869 163179 221897
rect 163207 221869 163241 221897
rect 163269 221869 178539 221897
rect 178567 221869 178601 221897
rect 178629 221869 193899 221897
rect 193927 221869 193961 221897
rect 193989 221869 209259 221897
rect 209287 221869 209321 221897
rect 209349 221869 224619 221897
rect 224647 221869 224681 221897
rect 224709 221869 239979 221897
rect 240007 221869 240041 221897
rect 240069 221869 256437 221897
rect 256465 221869 256499 221897
rect 256527 221869 256561 221897
rect 256589 221869 256623 221897
rect 256651 221869 265437 221897
rect 265465 221869 265499 221897
rect 265527 221869 265561 221897
rect 265589 221869 265623 221897
rect 265651 221869 274437 221897
rect 274465 221869 274499 221897
rect 274527 221869 274561 221897
rect 274589 221869 274623 221897
rect 274651 221869 283437 221897
rect 283465 221869 283499 221897
rect 283527 221869 283561 221897
rect 283589 221869 283623 221897
rect 283651 221869 292437 221897
rect 292465 221869 292499 221897
rect 292527 221869 292561 221897
rect 292589 221869 292623 221897
rect 292651 221869 299736 221897
rect 299764 221869 299798 221897
rect 299826 221869 299860 221897
rect 299888 221869 299922 221897
rect 299950 221869 299998 221897
rect -6 221835 299998 221869
rect -6 221807 42 221835
rect 70 221807 104 221835
rect 132 221807 166 221835
rect 194 221807 228 221835
rect 256 221807 4437 221835
rect 4465 221807 4499 221835
rect 4527 221807 4561 221835
rect 4589 221807 4623 221835
rect 4651 221807 13437 221835
rect 13465 221807 13499 221835
rect 13527 221807 13561 221835
rect 13589 221807 13623 221835
rect 13651 221807 22437 221835
rect 22465 221807 22499 221835
rect 22527 221807 22561 221835
rect 22589 221807 22623 221835
rect 22651 221807 24939 221835
rect 24967 221807 25001 221835
rect 25029 221807 31437 221835
rect 31465 221807 31499 221835
rect 31527 221807 31561 221835
rect 31589 221807 31623 221835
rect 31651 221807 40299 221835
rect 40327 221807 40361 221835
rect 40389 221807 55659 221835
rect 55687 221807 55721 221835
rect 55749 221807 71019 221835
rect 71047 221807 71081 221835
rect 71109 221807 86379 221835
rect 86407 221807 86441 221835
rect 86469 221807 101739 221835
rect 101767 221807 101801 221835
rect 101829 221807 117099 221835
rect 117127 221807 117161 221835
rect 117189 221807 132459 221835
rect 132487 221807 132521 221835
rect 132549 221807 147819 221835
rect 147847 221807 147881 221835
rect 147909 221807 163179 221835
rect 163207 221807 163241 221835
rect 163269 221807 178539 221835
rect 178567 221807 178601 221835
rect 178629 221807 193899 221835
rect 193927 221807 193961 221835
rect 193989 221807 209259 221835
rect 209287 221807 209321 221835
rect 209349 221807 224619 221835
rect 224647 221807 224681 221835
rect 224709 221807 239979 221835
rect 240007 221807 240041 221835
rect 240069 221807 256437 221835
rect 256465 221807 256499 221835
rect 256527 221807 256561 221835
rect 256589 221807 256623 221835
rect 256651 221807 265437 221835
rect 265465 221807 265499 221835
rect 265527 221807 265561 221835
rect 265589 221807 265623 221835
rect 265651 221807 274437 221835
rect 274465 221807 274499 221835
rect 274527 221807 274561 221835
rect 274589 221807 274623 221835
rect 274651 221807 283437 221835
rect 283465 221807 283499 221835
rect 283527 221807 283561 221835
rect 283589 221807 283623 221835
rect 283651 221807 292437 221835
rect 292465 221807 292499 221835
rect 292527 221807 292561 221835
rect 292589 221807 292623 221835
rect 292651 221807 299736 221835
rect 299764 221807 299798 221835
rect 299826 221807 299860 221835
rect 299888 221807 299922 221835
rect 299950 221807 299998 221835
rect -6 221773 299998 221807
rect -6 221745 42 221773
rect 70 221745 104 221773
rect 132 221745 166 221773
rect 194 221745 228 221773
rect 256 221745 4437 221773
rect 4465 221745 4499 221773
rect 4527 221745 4561 221773
rect 4589 221745 4623 221773
rect 4651 221745 13437 221773
rect 13465 221745 13499 221773
rect 13527 221745 13561 221773
rect 13589 221745 13623 221773
rect 13651 221745 22437 221773
rect 22465 221745 22499 221773
rect 22527 221745 22561 221773
rect 22589 221745 22623 221773
rect 22651 221745 24939 221773
rect 24967 221745 25001 221773
rect 25029 221745 31437 221773
rect 31465 221745 31499 221773
rect 31527 221745 31561 221773
rect 31589 221745 31623 221773
rect 31651 221745 40299 221773
rect 40327 221745 40361 221773
rect 40389 221745 55659 221773
rect 55687 221745 55721 221773
rect 55749 221745 71019 221773
rect 71047 221745 71081 221773
rect 71109 221745 86379 221773
rect 86407 221745 86441 221773
rect 86469 221745 101739 221773
rect 101767 221745 101801 221773
rect 101829 221745 117099 221773
rect 117127 221745 117161 221773
rect 117189 221745 132459 221773
rect 132487 221745 132521 221773
rect 132549 221745 147819 221773
rect 147847 221745 147881 221773
rect 147909 221745 163179 221773
rect 163207 221745 163241 221773
rect 163269 221745 178539 221773
rect 178567 221745 178601 221773
rect 178629 221745 193899 221773
rect 193927 221745 193961 221773
rect 193989 221745 209259 221773
rect 209287 221745 209321 221773
rect 209349 221745 224619 221773
rect 224647 221745 224681 221773
rect 224709 221745 239979 221773
rect 240007 221745 240041 221773
rect 240069 221745 256437 221773
rect 256465 221745 256499 221773
rect 256527 221745 256561 221773
rect 256589 221745 256623 221773
rect 256651 221745 265437 221773
rect 265465 221745 265499 221773
rect 265527 221745 265561 221773
rect 265589 221745 265623 221773
rect 265651 221745 274437 221773
rect 274465 221745 274499 221773
rect 274527 221745 274561 221773
rect 274589 221745 274623 221773
rect 274651 221745 283437 221773
rect 283465 221745 283499 221773
rect 283527 221745 283561 221773
rect 283589 221745 283623 221773
rect 283651 221745 292437 221773
rect 292465 221745 292499 221773
rect 292527 221745 292561 221773
rect 292589 221745 292623 221773
rect 292651 221745 299736 221773
rect 299764 221745 299798 221773
rect 299826 221745 299860 221773
rect 299888 221745 299922 221773
rect 299950 221745 299998 221773
rect -6 221697 299998 221745
rect -6 218959 299998 219007
rect -6 218931 522 218959
rect 550 218931 584 218959
rect 612 218931 646 218959
rect 674 218931 708 218959
rect 736 218931 2577 218959
rect 2605 218931 2639 218959
rect 2667 218931 2701 218959
rect 2729 218931 2763 218959
rect 2791 218931 11577 218959
rect 11605 218931 11639 218959
rect 11667 218931 11701 218959
rect 11729 218931 11763 218959
rect 11791 218931 17259 218959
rect 17287 218931 17321 218959
rect 17349 218931 20577 218959
rect 20605 218931 20639 218959
rect 20667 218931 20701 218959
rect 20729 218931 20763 218959
rect 20791 218931 29577 218959
rect 29605 218931 29639 218959
rect 29667 218931 29701 218959
rect 29729 218931 29763 218959
rect 29791 218931 32619 218959
rect 32647 218931 32681 218959
rect 32709 218931 47979 218959
rect 48007 218931 48041 218959
rect 48069 218931 63339 218959
rect 63367 218931 63401 218959
rect 63429 218931 78699 218959
rect 78727 218931 78761 218959
rect 78789 218931 94059 218959
rect 94087 218931 94121 218959
rect 94149 218931 109419 218959
rect 109447 218931 109481 218959
rect 109509 218931 124779 218959
rect 124807 218931 124841 218959
rect 124869 218931 140139 218959
rect 140167 218931 140201 218959
rect 140229 218931 155499 218959
rect 155527 218931 155561 218959
rect 155589 218931 170859 218959
rect 170887 218931 170921 218959
rect 170949 218931 186219 218959
rect 186247 218931 186281 218959
rect 186309 218931 201579 218959
rect 201607 218931 201641 218959
rect 201669 218931 216939 218959
rect 216967 218931 217001 218959
rect 217029 218931 232299 218959
rect 232327 218931 232361 218959
rect 232389 218931 247659 218959
rect 247687 218931 247721 218959
rect 247749 218931 254577 218959
rect 254605 218931 254639 218959
rect 254667 218931 254701 218959
rect 254729 218931 254763 218959
rect 254791 218931 263577 218959
rect 263605 218931 263639 218959
rect 263667 218931 263701 218959
rect 263729 218931 263763 218959
rect 263791 218931 272577 218959
rect 272605 218931 272639 218959
rect 272667 218931 272701 218959
rect 272729 218931 272763 218959
rect 272791 218931 281577 218959
rect 281605 218931 281639 218959
rect 281667 218931 281701 218959
rect 281729 218931 281763 218959
rect 281791 218931 290577 218959
rect 290605 218931 290639 218959
rect 290667 218931 290701 218959
rect 290729 218931 290763 218959
rect 290791 218931 299256 218959
rect 299284 218931 299318 218959
rect 299346 218931 299380 218959
rect 299408 218931 299442 218959
rect 299470 218931 299998 218959
rect -6 218897 299998 218931
rect -6 218869 522 218897
rect 550 218869 584 218897
rect 612 218869 646 218897
rect 674 218869 708 218897
rect 736 218869 2577 218897
rect 2605 218869 2639 218897
rect 2667 218869 2701 218897
rect 2729 218869 2763 218897
rect 2791 218869 11577 218897
rect 11605 218869 11639 218897
rect 11667 218869 11701 218897
rect 11729 218869 11763 218897
rect 11791 218869 17259 218897
rect 17287 218869 17321 218897
rect 17349 218869 20577 218897
rect 20605 218869 20639 218897
rect 20667 218869 20701 218897
rect 20729 218869 20763 218897
rect 20791 218869 29577 218897
rect 29605 218869 29639 218897
rect 29667 218869 29701 218897
rect 29729 218869 29763 218897
rect 29791 218869 32619 218897
rect 32647 218869 32681 218897
rect 32709 218869 47979 218897
rect 48007 218869 48041 218897
rect 48069 218869 63339 218897
rect 63367 218869 63401 218897
rect 63429 218869 78699 218897
rect 78727 218869 78761 218897
rect 78789 218869 94059 218897
rect 94087 218869 94121 218897
rect 94149 218869 109419 218897
rect 109447 218869 109481 218897
rect 109509 218869 124779 218897
rect 124807 218869 124841 218897
rect 124869 218869 140139 218897
rect 140167 218869 140201 218897
rect 140229 218869 155499 218897
rect 155527 218869 155561 218897
rect 155589 218869 170859 218897
rect 170887 218869 170921 218897
rect 170949 218869 186219 218897
rect 186247 218869 186281 218897
rect 186309 218869 201579 218897
rect 201607 218869 201641 218897
rect 201669 218869 216939 218897
rect 216967 218869 217001 218897
rect 217029 218869 232299 218897
rect 232327 218869 232361 218897
rect 232389 218869 247659 218897
rect 247687 218869 247721 218897
rect 247749 218869 254577 218897
rect 254605 218869 254639 218897
rect 254667 218869 254701 218897
rect 254729 218869 254763 218897
rect 254791 218869 263577 218897
rect 263605 218869 263639 218897
rect 263667 218869 263701 218897
rect 263729 218869 263763 218897
rect 263791 218869 272577 218897
rect 272605 218869 272639 218897
rect 272667 218869 272701 218897
rect 272729 218869 272763 218897
rect 272791 218869 281577 218897
rect 281605 218869 281639 218897
rect 281667 218869 281701 218897
rect 281729 218869 281763 218897
rect 281791 218869 290577 218897
rect 290605 218869 290639 218897
rect 290667 218869 290701 218897
rect 290729 218869 290763 218897
rect 290791 218869 299256 218897
rect 299284 218869 299318 218897
rect 299346 218869 299380 218897
rect 299408 218869 299442 218897
rect 299470 218869 299998 218897
rect -6 218835 299998 218869
rect -6 218807 522 218835
rect 550 218807 584 218835
rect 612 218807 646 218835
rect 674 218807 708 218835
rect 736 218807 2577 218835
rect 2605 218807 2639 218835
rect 2667 218807 2701 218835
rect 2729 218807 2763 218835
rect 2791 218807 11577 218835
rect 11605 218807 11639 218835
rect 11667 218807 11701 218835
rect 11729 218807 11763 218835
rect 11791 218807 17259 218835
rect 17287 218807 17321 218835
rect 17349 218807 20577 218835
rect 20605 218807 20639 218835
rect 20667 218807 20701 218835
rect 20729 218807 20763 218835
rect 20791 218807 29577 218835
rect 29605 218807 29639 218835
rect 29667 218807 29701 218835
rect 29729 218807 29763 218835
rect 29791 218807 32619 218835
rect 32647 218807 32681 218835
rect 32709 218807 47979 218835
rect 48007 218807 48041 218835
rect 48069 218807 63339 218835
rect 63367 218807 63401 218835
rect 63429 218807 78699 218835
rect 78727 218807 78761 218835
rect 78789 218807 94059 218835
rect 94087 218807 94121 218835
rect 94149 218807 109419 218835
rect 109447 218807 109481 218835
rect 109509 218807 124779 218835
rect 124807 218807 124841 218835
rect 124869 218807 140139 218835
rect 140167 218807 140201 218835
rect 140229 218807 155499 218835
rect 155527 218807 155561 218835
rect 155589 218807 170859 218835
rect 170887 218807 170921 218835
rect 170949 218807 186219 218835
rect 186247 218807 186281 218835
rect 186309 218807 201579 218835
rect 201607 218807 201641 218835
rect 201669 218807 216939 218835
rect 216967 218807 217001 218835
rect 217029 218807 232299 218835
rect 232327 218807 232361 218835
rect 232389 218807 247659 218835
rect 247687 218807 247721 218835
rect 247749 218807 254577 218835
rect 254605 218807 254639 218835
rect 254667 218807 254701 218835
rect 254729 218807 254763 218835
rect 254791 218807 263577 218835
rect 263605 218807 263639 218835
rect 263667 218807 263701 218835
rect 263729 218807 263763 218835
rect 263791 218807 272577 218835
rect 272605 218807 272639 218835
rect 272667 218807 272701 218835
rect 272729 218807 272763 218835
rect 272791 218807 281577 218835
rect 281605 218807 281639 218835
rect 281667 218807 281701 218835
rect 281729 218807 281763 218835
rect 281791 218807 290577 218835
rect 290605 218807 290639 218835
rect 290667 218807 290701 218835
rect 290729 218807 290763 218835
rect 290791 218807 299256 218835
rect 299284 218807 299318 218835
rect 299346 218807 299380 218835
rect 299408 218807 299442 218835
rect 299470 218807 299998 218835
rect -6 218773 299998 218807
rect -6 218745 522 218773
rect 550 218745 584 218773
rect 612 218745 646 218773
rect 674 218745 708 218773
rect 736 218745 2577 218773
rect 2605 218745 2639 218773
rect 2667 218745 2701 218773
rect 2729 218745 2763 218773
rect 2791 218745 11577 218773
rect 11605 218745 11639 218773
rect 11667 218745 11701 218773
rect 11729 218745 11763 218773
rect 11791 218745 17259 218773
rect 17287 218745 17321 218773
rect 17349 218745 20577 218773
rect 20605 218745 20639 218773
rect 20667 218745 20701 218773
rect 20729 218745 20763 218773
rect 20791 218745 29577 218773
rect 29605 218745 29639 218773
rect 29667 218745 29701 218773
rect 29729 218745 29763 218773
rect 29791 218745 32619 218773
rect 32647 218745 32681 218773
rect 32709 218745 47979 218773
rect 48007 218745 48041 218773
rect 48069 218745 63339 218773
rect 63367 218745 63401 218773
rect 63429 218745 78699 218773
rect 78727 218745 78761 218773
rect 78789 218745 94059 218773
rect 94087 218745 94121 218773
rect 94149 218745 109419 218773
rect 109447 218745 109481 218773
rect 109509 218745 124779 218773
rect 124807 218745 124841 218773
rect 124869 218745 140139 218773
rect 140167 218745 140201 218773
rect 140229 218745 155499 218773
rect 155527 218745 155561 218773
rect 155589 218745 170859 218773
rect 170887 218745 170921 218773
rect 170949 218745 186219 218773
rect 186247 218745 186281 218773
rect 186309 218745 201579 218773
rect 201607 218745 201641 218773
rect 201669 218745 216939 218773
rect 216967 218745 217001 218773
rect 217029 218745 232299 218773
rect 232327 218745 232361 218773
rect 232389 218745 247659 218773
rect 247687 218745 247721 218773
rect 247749 218745 254577 218773
rect 254605 218745 254639 218773
rect 254667 218745 254701 218773
rect 254729 218745 254763 218773
rect 254791 218745 263577 218773
rect 263605 218745 263639 218773
rect 263667 218745 263701 218773
rect 263729 218745 263763 218773
rect 263791 218745 272577 218773
rect 272605 218745 272639 218773
rect 272667 218745 272701 218773
rect 272729 218745 272763 218773
rect 272791 218745 281577 218773
rect 281605 218745 281639 218773
rect 281667 218745 281701 218773
rect 281729 218745 281763 218773
rect 281791 218745 290577 218773
rect 290605 218745 290639 218773
rect 290667 218745 290701 218773
rect 290729 218745 290763 218773
rect 290791 218745 299256 218773
rect 299284 218745 299318 218773
rect 299346 218745 299380 218773
rect 299408 218745 299442 218773
rect 299470 218745 299998 218773
rect -6 218697 299998 218745
rect -6 212959 299998 213007
rect -6 212931 42 212959
rect 70 212931 104 212959
rect 132 212931 166 212959
rect 194 212931 228 212959
rect 256 212931 4437 212959
rect 4465 212931 4499 212959
rect 4527 212931 4561 212959
rect 4589 212931 4623 212959
rect 4651 212931 13437 212959
rect 13465 212931 13499 212959
rect 13527 212931 13561 212959
rect 13589 212931 13623 212959
rect 13651 212931 22437 212959
rect 22465 212931 22499 212959
rect 22527 212931 22561 212959
rect 22589 212931 22623 212959
rect 22651 212931 24939 212959
rect 24967 212931 25001 212959
rect 25029 212931 31437 212959
rect 31465 212931 31499 212959
rect 31527 212931 31561 212959
rect 31589 212931 31623 212959
rect 31651 212931 40299 212959
rect 40327 212931 40361 212959
rect 40389 212931 55659 212959
rect 55687 212931 55721 212959
rect 55749 212931 71019 212959
rect 71047 212931 71081 212959
rect 71109 212931 86379 212959
rect 86407 212931 86441 212959
rect 86469 212931 101739 212959
rect 101767 212931 101801 212959
rect 101829 212931 117099 212959
rect 117127 212931 117161 212959
rect 117189 212931 132459 212959
rect 132487 212931 132521 212959
rect 132549 212931 147819 212959
rect 147847 212931 147881 212959
rect 147909 212931 163179 212959
rect 163207 212931 163241 212959
rect 163269 212931 178539 212959
rect 178567 212931 178601 212959
rect 178629 212931 193899 212959
rect 193927 212931 193961 212959
rect 193989 212931 209259 212959
rect 209287 212931 209321 212959
rect 209349 212931 224619 212959
rect 224647 212931 224681 212959
rect 224709 212931 239979 212959
rect 240007 212931 240041 212959
rect 240069 212931 256437 212959
rect 256465 212931 256499 212959
rect 256527 212931 256561 212959
rect 256589 212931 256623 212959
rect 256651 212931 265437 212959
rect 265465 212931 265499 212959
rect 265527 212931 265561 212959
rect 265589 212931 265623 212959
rect 265651 212931 274437 212959
rect 274465 212931 274499 212959
rect 274527 212931 274561 212959
rect 274589 212931 274623 212959
rect 274651 212931 283437 212959
rect 283465 212931 283499 212959
rect 283527 212931 283561 212959
rect 283589 212931 283623 212959
rect 283651 212931 292437 212959
rect 292465 212931 292499 212959
rect 292527 212931 292561 212959
rect 292589 212931 292623 212959
rect 292651 212931 299736 212959
rect 299764 212931 299798 212959
rect 299826 212931 299860 212959
rect 299888 212931 299922 212959
rect 299950 212931 299998 212959
rect -6 212897 299998 212931
rect -6 212869 42 212897
rect 70 212869 104 212897
rect 132 212869 166 212897
rect 194 212869 228 212897
rect 256 212869 4437 212897
rect 4465 212869 4499 212897
rect 4527 212869 4561 212897
rect 4589 212869 4623 212897
rect 4651 212869 13437 212897
rect 13465 212869 13499 212897
rect 13527 212869 13561 212897
rect 13589 212869 13623 212897
rect 13651 212869 22437 212897
rect 22465 212869 22499 212897
rect 22527 212869 22561 212897
rect 22589 212869 22623 212897
rect 22651 212869 24939 212897
rect 24967 212869 25001 212897
rect 25029 212869 31437 212897
rect 31465 212869 31499 212897
rect 31527 212869 31561 212897
rect 31589 212869 31623 212897
rect 31651 212869 40299 212897
rect 40327 212869 40361 212897
rect 40389 212869 55659 212897
rect 55687 212869 55721 212897
rect 55749 212869 71019 212897
rect 71047 212869 71081 212897
rect 71109 212869 86379 212897
rect 86407 212869 86441 212897
rect 86469 212869 101739 212897
rect 101767 212869 101801 212897
rect 101829 212869 117099 212897
rect 117127 212869 117161 212897
rect 117189 212869 132459 212897
rect 132487 212869 132521 212897
rect 132549 212869 147819 212897
rect 147847 212869 147881 212897
rect 147909 212869 163179 212897
rect 163207 212869 163241 212897
rect 163269 212869 178539 212897
rect 178567 212869 178601 212897
rect 178629 212869 193899 212897
rect 193927 212869 193961 212897
rect 193989 212869 209259 212897
rect 209287 212869 209321 212897
rect 209349 212869 224619 212897
rect 224647 212869 224681 212897
rect 224709 212869 239979 212897
rect 240007 212869 240041 212897
rect 240069 212869 256437 212897
rect 256465 212869 256499 212897
rect 256527 212869 256561 212897
rect 256589 212869 256623 212897
rect 256651 212869 265437 212897
rect 265465 212869 265499 212897
rect 265527 212869 265561 212897
rect 265589 212869 265623 212897
rect 265651 212869 274437 212897
rect 274465 212869 274499 212897
rect 274527 212869 274561 212897
rect 274589 212869 274623 212897
rect 274651 212869 283437 212897
rect 283465 212869 283499 212897
rect 283527 212869 283561 212897
rect 283589 212869 283623 212897
rect 283651 212869 292437 212897
rect 292465 212869 292499 212897
rect 292527 212869 292561 212897
rect 292589 212869 292623 212897
rect 292651 212869 299736 212897
rect 299764 212869 299798 212897
rect 299826 212869 299860 212897
rect 299888 212869 299922 212897
rect 299950 212869 299998 212897
rect -6 212835 299998 212869
rect -6 212807 42 212835
rect 70 212807 104 212835
rect 132 212807 166 212835
rect 194 212807 228 212835
rect 256 212807 4437 212835
rect 4465 212807 4499 212835
rect 4527 212807 4561 212835
rect 4589 212807 4623 212835
rect 4651 212807 13437 212835
rect 13465 212807 13499 212835
rect 13527 212807 13561 212835
rect 13589 212807 13623 212835
rect 13651 212807 22437 212835
rect 22465 212807 22499 212835
rect 22527 212807 22561 212835
rect 22589 212807 22623 212835
rect 22651 212807 24939 212835
rect 24967 212807 25001 212835
rect 25029 212807 31437 212835
rect 31465 212807 31499 212835
rect 31527 212807 31561 212835
rect 31589 212807 31623 212835
rect 31651 212807 40299 212835
rect 40327 212807 40361 212835
rect 40389 212807 55659 212835
rect 55687 212807 55721 212835
rect 55749 212807 71019 212835
rect 71047 212807 71081 212835
rect 71109 212807 86379 212835
rect 86407 212807 86441 212835
rect 86469 212807 101739 212835
rect 101767 212807 101801 212835
rect 101829 212807 117099 212835
rect 117127 212807 117161 212835
rect 117189 212807 132459 212835
rect 132487 212807 132521 212835
rect 132549 212807 147819 212835
rect 147847 212807 147881 212835
rect 147909 212807 163179 212835
rect 163207 212807 163241 212835
rect 163269 212807 178539 212835
rect 178567 212807 178601 212835
rect 178629 212807 193899 212835
rect 193927 212807 193961 212835
rect 193989 212807 209259 212835
rect 209287 212807 209321 212835
rect 209349 212807 224619 212835
rect 224647 212807 224681 212835
rect 224709 212807 239979 212835
rect 240007 212807 240041 212835
rect 240069 212807 256437 212835
rect 256465 212807 256499 212835
rect 256527 212807 256561 212835
rect 256589 212807 256623 212835
rect 256651 212807 265437 212835
rect 265465 212807 265499 212835
rect 265527 212807 265561 212835
rect 265589 212807 265623 212835
rect 265651 212807 274437 212835
rect 274465 212807 274499 212835
rect 274527 212807 274561 212835
rect 274589 212807 274623 212835
rect 274651 212807 283437 212835
rect 283465 212807 283499 212835
rect 283527 212807 283561 212835
rect 283589 212807 283623 212835
rect 283651 212807 292437 212835
rect 292465 212807 292499 212835
rect 292527 212807 292561 212835
rect 292589 212807 292623 212835
rect 292651 212807 299736 212835
rect 299764 212807 299798 212835
rect 299826 212807 299860 212835
rect 299888 212807 299922 212835
rect 299950 212807 299998 212835
rect -6 212773 299998 212807
rect -6 212745 42 212773
rect 70 212745 104 212773
rect 132 212745 166 212773
rect 194 212745 228 212773
rect 256 212745 4437 212773
rect 4465 212745 4499 212773
rect 4527 212745 4561 212773
rect 4589 212745 4623 212773
rect 4651 212745 13437 212773
rect 13465 212745 13499 212773
rect 13527 212745 13561 212773
rect 13589 212745 13623 212773
rect 13651 212745 22437 212773
rect 22465 212745 22499 212773
rect 22527 212745 22561 212773
rect 22589 212745 22623 212773
rect 22651 212745 24939 212773
rect 24967 212745 25001 212773
rect 25029 212745 31437 212773
rect 31465 212745 31499 212773
rect 31527 212745 31561 212773
rect 31589 212745 31623 212773
rect 31651 212745 40299 212773
rect 40327 212745 40361 212773
rect 40389 212745 55659 212773
rect 55687 212745 55721 212773
rect 55749 212745 71019 212773
rect 71047 212745 71081 212773
rect 71109 212745 86379 212773
rect 86407 212745 86441 212773
rect 86469 212745 101739 212773
rect 101767 212745 101801 212773
rect 101829 212745 117099 212773
rect 117127 212745 117161 212773
rect 117189 212745 132459 212773
rect 132487 212745 132521 212773
rect 132549 212745 147819 212773
rect 147847 212745 147881 212773
rect 147909 212745 163179 212773
rect 163207 212745 163241 212773
rect 163269 212745 178539 212773
rect 178567 212745 178601 212773
rect 178629 212745 193899 212773
rect 193927 212745 193961 212773
rect 193989 212745 209259 212773
rect 209287 212745 209321 212773
rect 209349 212745 224619 212773
rect 224647 212745 224681 212773
rect 224709 212745 239979 212773
rect 240007 212745 240041 212773
rect 240069 212745 256437 212773
rect 256465 212745 256499 212773
rect 256527 212745 256561 212773
rect 256589 212745 256623 212773
rect 256651 212745 265437 212773
rect 265465 212745 265499 212773
rect 265527 212745 265561 212773
rect 265589 212745 265623 212773
rect 265651 212745 274437 212773
rect 274465 212745 274499 212773
rect 274527 212745 274561 212773
rect 274589 212745 274623 212773
rect 274651 212745 283437 212773
rect 283465 212745 283499 212773
rect 283527 212745 283561 212773
rect 283589 212745 283623 212773
rect 283651 212745 292437 212773
rect 292465 212745 292499 212773
rect 292527 212745 292561 212773
rect 292589 212745 292623 212773
rect 292651 212745 299736 212773
rect 299764 212745 299798 212773
rect 299826 212745 299860 212773
rect 299888 212745 299922 212773
rect 299950 212745 299998 212773
rect -6 212697 299998 212745
rect -6 209959 299998 210007
rect -6 209931 522 209959
rect 550 209931 584 209959
rect 612 209931 646 209959
rect 674 209931 708 209959
rect 736 209931 2577 209959
rect 2605 209931 2639 209959
rect 2667 209931 2701 209959
rect 2729 209931 2763 209959
rect 2791 209931 11577 209959
rect 11605 209931 11639 209959
rect 11667 209931 11701 209959
rect 11729 209931 11763 209959
rect 11791 209931 17259 209959
rect 17287 209931 17321 209959
rect 17349 209931 20577 209959
rect 20605 209931 20639 209959
rect 20667 209931 20701 209959
rect 20729 209931 20763 209959
rect 20791 209931 29577 209959
rect 29605 209931 29639 209959
rect 29667 209931 29701 209959
rect 29729 209931 29763 209959
rect 29791 209931 32619 209959
rect 32647 209931 32681 209959
rect 32709 209931 47979 209959
rect 48007 209931 48041 209959
rect 48069 209931 63339 209959
rect 63367 209931 63401 209959
rect 63429 209931 78699 209959
rect 78727 209931 78761 209959
rect 78789 209931 94059 209959
rect 94087 209931 94121 209959
rect 94149 209931 109419 209959
rect 109447 209931 109481 209959
rect 109509 209931 124779 209959
rect 124807 209931 124841 209959
rect 124869 209931 140139 209959
rect 140167 209931 140201 209959
rect 140229 209931 155499 209959
rect 155527 209931 155561 209959
rect 155589 209931 170859 209959
rect 170887 209931 170921 209959
rect 170949 209931 186219 209959
rect 186247 209931 186281 209959
rect 186309 209931 201579 209959
rect 201607 209931 201641 209959
rect 201669 209931 216939 209959
rect 216967 209931 217001 209959
rect 217029 209931 232299 209959
rect 232327 209931 232361 209959
rect 232389 209931 247659 209959
rect 247687 209931 247721 209959
rect 247749 209931 254577 209959
rect 254605 209931 254639 209959
rect 254667 209931 254701 209959
rect 254729 209931 254763 209959
rect 254791 209931 263577 209959
rect 263605 209931 263639 209959
rect 263667 209931 263701 209959
rect 263729 209931 263763 209959
rect 263791 209931 272577 209959
rect 272605 209931 272639 209959
rect 272667 209931 272701 209959
rect 272729 209931 272763 209959
rect 272791 209931 281577 209959
rect 281605 209931 281639 209959
rect 281667 209931 281701 209959
rect 281729 209931 281763 209959
rect 281791 209931 290577 209959
rect 290605 209931 290639 209959
rect 290667 209931 290701 209959
rect 290729 209931 290763 209959
rect 290791 209931 299256 209959
rect 299284 209931 299318 209959
rect 299346 209931 299380 209959
rect 299408 209931 299442 209959
rect 299470 209931 299998 209959
rect -6 209897 299998 209931
rect -6 209869 522 209897
rect 550 209869 584 209897
rect 612 209869 646 209897
rect 674 209869 708 209897
rect 736 209869 2577 209897
rect 2605 209869 2639 209897
rect 2667 209869 2701 209897
rect 2729 209869 2763 209897
rect 2791 209869 11577 209897
rect 11605 209869 11639 209897
rect 11667 209869 11701 209897
rect 11729 209869 11763 209897
rect 11791 209869 17259 209897
rect 17287 209869 17321 209897
rect 17349 209869 20577 209897
rect 20605 209869 20639 209897
rect 20667 209869 20701 209897
rect 20729 209869 20763 209897
rect 20791 209869 29577 209897
rect 29605 209869 29639 209897
rect 29667 209869 29701 209897
rect 29729 209869 29763 209897
rect 29791 209869 32619 209897
rect 32647 209869 32681 209897
rect 32709 209869 47979 209897
rect 48007 209869 48041 209897
rect 48069 209869 63339 209897
rect 63367 209869 63401 209897
rect 63429 209869 78699 209897
rect 78727 209869 78761 209897
rect 78789 209869 94059 209897
rect 94087 209869 94121 209897
rect 94149 209869 109419 209897
rect 109447 209869 109481 209897
rect 109509 209869 124779 209897
rect 124807 209869 124841 209897
rect 124869 209869 140139 209897
rect 140167 209869 140201 209897
rect 140229 209869 155499 209897
rect 155527 209869 155561 209897
rect 155589 209869 170859 209897
rect 170887 209869 170921 209897
rect 170949 209869 186219 209897
rect 186247 209869 186281 209897
rect 186309 209869 201579 209897
rect 201607 209869 201641 209897
rect 201669 209869 216939 209897
rect 216967 209869 217001 209897
rect 217029 209869 232299 209897
rect 232327 209869 232361 209897
rect 232389 209869 247659 209897
rect 247687 209869 247721 209897
rect 247749 209869 254577 209897
rect 254605 209869 254639 209897
rect 254667 209869 254701 209897
rect 254729 209869 254763 209897
rect 254791 209869 263577 209897
rect 263605 209869 263639 209897
rect 263667 209869 263701 209897
rect 263729 209869 263763 209897
rect 263791 209869 272577 209897
rect 272605 209869 272639 209897
rect 272667 209869 272701 209897
rect 272729 209869 272763 209897
rect 272791 209869 281577 209897
rect 281605 209869 281639 209897
rect 281667 209869 281701 209897
rect 281729 209869 281763 209897
rect 281791 209869 290577 209897
rect 290605 209869 290639 209897
rect 290667 209869 290701 209897
rect 290729 209869 290763 209897
rect 290791 209869 299256 209897
rect 299284 209869 299318 209897
rect 299346 209869 299380 209897
rect 299408 209869 299442 209897
rect 299470 209869 299998 209897
rect -6 209835 299998 209869
rect -6 209807 522 209835
rect 550 209807 584 209835
rect 612 209807 646 209835
rect 674 209807 708 209835
rect 736 209807 2577 209835
rect 2605 209807 2639 209835
rect 2667 209807 2701 209835
rect 2729 209807 2763 209835
rect 2791 209807 11577 209835
rect 11605 209807 11639 209835
rect 11667 209807 11701 209835
rect 11729 209807 11763 209835
rect 11791 209807 17259 209835
rect 17287 209807 17321 209835
rect 17349 209807 20577 209835
rect 20605 209807 20639 209835
rect 20667 209807 20701 209835
rect 20729 209807 20763 209835
rect 20791 209807 29577 209835
rect 29605 209807 29639 209835
rect 29667 209807 29701 209835
rect 29729 209807 29763 209835
rect 29791 209807 32619 209835
rect 32647 209807 32681 209835
rect 32709 209807 47979 209835
rect 48007 209807 48041 209835
rect 48069 209807 63339 209835
rect 63367 209807 63401 209835
rect 63429 209807 78699 209835
rect 78727 209807 78761 209835
rect 78789 209807 94059 209835
rect 94087 209807 94121 209835
rect 94149 209807 109419 209835
rect 109447 209807 109481 209835
rect 109509 209807 124779 209835
rect 124807 209807 124841 209835
rect 124869 209807 140139 209835
rect 140167 209807 140201 209835
rect 140229 209807 155499 209835
rect 155527 209807 155561 209835
rect 155589 209807 170859 209835
rect 170887 209807 170921 209835
rect 170949 209807 186219 209835
rect 186247 209807 186281 209835
rect 186309 209807 201579 209835
rect 201607 209807 201641 209835
rect 201669 209807 216939 209835
rect 216967 209807 217001 209835
rect 217029 209807 232299 209835
rect 232327 209807 232361 209835
rect 232389 209807 247659 209835
rect 247687 209807 247721 209835
rect 247749 209807 254577 209835
rect 254605 209807 254639 209835
rect 254667 209807 254701 209835
rect 254729 209807 254763 209835
rect 254791 209807 263577 209835
rect 263605 209807 263639 209835
rect 263667 209807 263701 209835
rect 263729 209807 263763 209835
rect 263791 209807 272577 209835
rect 272605 209807 272639 209835
rect 272667 209807 272701 209835
rect 272729 209807 272763 209835
rect 272791 209807 281577 209835
rect 281605 209807 281639 209835
rect 281667 209807 281701 209835
rect 281729 209807 281763 209835
rect 281791 209807 290577 209835
rect 290605 209807 290639 209835
rect 290667 209807 290701 209835
rect 290729 209807 290763 209835
rect 290791 209807 299256 209835
rect 299284 209807 299318 209835
rect 299346 209807 299380 209835
rect 299408 209807 299442 209835
rect 299470 209807 299998 209835
rect -6 209773 299998 209807
rect -6 209745 522 209773
rect 550 209745 584 209773
rect 612 209745 646 209773
rect 674 209745 708 209773
rect 736 209745 2577 209773
rect 2605 209745 2639 209773
rect 2667 209745 2701 209773
rect 2729 209745 2763 209773
rect 2791 209745 11577 209773
rect 11605 209745 11639 209773
rect 11667 209745 11701 209773
rect 11729 209745 11763 209773
rect 11791 209745 17259 209773
rect 17287 209745 17321 209773
rect 17349 209745 20577 209773
rect 20605 209745 20639 209773
rect 20667 209745 20701 209773
rect 20729 209745 20763 209773
rect 20791 209745 29577 209773
rect 29605 209745 29639 209773
rect 29667 209745 29701 209773
rect 29729 209745 29763 209773
rect 29791 209745 32619 209773
rect 32647 209745 32681 209773
rect 32709 209745 47979 209773
rect 48007 209745 48041 209773
rect 48069 209745 63339 209773
rect 63367 209745 63401 209773
rect 63429 209745 78699 209773
rect 78727 209745 78761 209773
rect 78789 209745 94059 209773
rect 94087 209745 94121 209773
rect 94149 209745 109419 209773
rect 109447 209745 109481 209773
rect 109509 209745 124779 209773
rect 124807 209745 124841 209773
rect 124869 209745 140139 209773
rect 140167 209745 140201 209773
rect 140229 209745 155499 209773
rect 155527 209745 155561 209773
rect 155589 209745 170859 209773
rect 170887 209745 170921 209773
rect 170949 209745 186219 209773
rect 186247 209745 186281 209773
rect 186309 209745 201579 209773
rect 201607 209745 201641 209773
rect 201669 209745 216939 209773
rect 216967 209745 217001 209773
rect 217029 209745 232299 209773
rect 232327 209745 232361 209773
rect 232389 209745 247659 209773
rect 247687 209745 247721 209773
rect 247749 209745 254577 209773
rect 254605 209745 254639 209773
rect 254667 209745 254701 209773
rect 254729 209745 254763 209773
rect 254791 209745 263577 209773
rect 263605 209745 263639 209773
rect 263667 209745 263701 209773
rect 263729 209745 263763 209773
rect 263791 209745 272577 209773
rect 272605 209745 272639 209773
rect 272667 209745 272701 209773
rect 272729 209745 272763 209773
rect 272791 209745 281577 209773
rect 281605 209745 281639 209773
rect 281667 209745 281701 209773
rect 281729 209745 281763 209773
rect 281791 209745 290577 209773
rect 290605 209745 290639 209773
rect 290667 209745 290701 209773
rect 290729 209745 290763 209773
rect 290791 209745 299256 209773
rect 299284 209745 299318 209773
rect 299346 209745 299380 209773
rect 299408 209745 299442 209773
rect 299470 209745 299998 209773
rect -6 209697 299998 209745
rect -6 203959 299998 204007
rect -6 203931 42 203959
rect 70 203931 104 203959
rect 132 203931 166 203959
rect 194 203931 228 203959
rect 256 203931 4437 203959
rect 4465 203931 4499 203959
rect 4527 203931 4561 203959
rect 4589 203931 4623 203959
rect 4651 203931 13437 203959
rect 13465 203931 13499 203959
rect 13527 203931 13561 203959
rect 13589 203931 13623 203959
rect 13651 203931 22437 203959
rect 22465 203931 22499 203959
rect 22527 203931 22561 203959
rect 22589 203931 22623 203959
rect 22651 203931 24939 203959
rect 24967 203931 25001 203959
rect 25029 203931 31437 203959
rect 31465 203931 31499 203959
rect 31527 203931 31561 203959
rect 31589 203931 31623 203959
rect 31651 203931 40299 203959
rect 40327 203931 40361 203959
rect 40389 203931 55659 203959
rect 55687 203931 55721 203959
rect 55749 203931 71019 203959
rect 71047 203931 71081 203959
rect 71109 203931 86379 203959
rect 86407 203931 86441 203959
rect 86469 203931 101739 203959
rect 101767 203931 101801 203959
rect 101829 203931 117099 203959
rect 117127 203931 117161 203959
rect 117189 203931 132459 203959
rect 132487 203931 132521 203959
rect 132549 203931 147819 203959
rect 147847 203931 147881 203959
rect 147909 203931 163179 203959
rect 163207 203931 163241 203959
rect 163269 203931 178539 203959
rect 178567 203931 178601 203959
rect 178629 203931 193899 203959
rect 193927 203931 193961 203959
rect 193989 203931 209259 203959
rect 209287 203931 209321 203959
rect 209349 203931 224619 203959
rect 224647 203931 224681 203959
rect 224709 203931 239979 203959
rect 240007 203931 240041 203959
rect 240069 203931 256437 203959
rect 256465 203931 256499 203959
rect 256527 203931 256561 203959
rect 256589 203931 256623 203959
rect 256651 203931 265437 203959
rect 265465 203931 265499 203959
rect 265527 203931 265561 203959
rect 265589 203931 265623 203959
rect 265651 203931 274437 203959
rect 274465 203931 274499 203959
rect 274527 203931 274561 203959
rect 274589 203931 274623 203959
rect 274651 203931 283437 203959
rect 283465 203931 283499 203959
rect 283527 203931 283561 203959
rect 283589 203931 283623 203959
rect 283651 203931 292437 203959
rect 292465 203931 292499 203959
rect 292527 203931 292561 203959
rect 292589 203931 292623 203959
rect 292651 203931 299736 203959
rect 299764 203931 299798 203959
rect 299826 203931 299860 203959
rect 299888 203931 299922 203959
rect 299950 203931 299998 203959
rect -6 203897 299998 203931
rect -6 203869 42 203897
rect 70 203869 104 203897
rect 132 203869 166 203897
rect 194 203869 228 203897
rect 256 203869 4437 203897
rect 4465 203869 4499 203897
rect 4527 203869 4561 203897
rect 4589 203869 4623 203897
rect 4651 203869 13437 203897
rect 13465 203869 13499 203897
rect 13527 203869 13561 203897
rect 13589 203869 13623 203897
rect 13651 203869 22437 203897
rect 22465 203869 22499 203897
rect 22527 203869 22561 203897
rect 22589 203869 22623 203897
rect 22651 203869 24939 203897
rect 24967 203869 25001 203897
rect 25029 203869 31437 203897
rect 31465 203869 31499 203897
rect 31527 203869 31561 203897
rect 31589 203869 31623 203897
rect 31651 203869 40299 203897
rect 40327 203869 40361 203897
rect 40389 203869 55659 203897
rect 55687 203869 55721 203897
rect 55749 203869 71019 203897
rect 71047 203869 71081 203897
rect 71109 203869 86379 203897
rect 86407 203869 86441 203897
rect 86469 203869 101739 203897
rect 101767 203869 101801 203897
rect 101829 203869 117099 203897
rect 117127 203869 117161 203897
rect 117189 203869 132459 203897
rect 132487 203869 132521 203897
rect 132549 203869 147819 203897
rect 147847 203869 147881 203897
rect 147909 203869 163179 203897
rect 163207 203869 163241 203897
rect 163269 203869 178539 203897
rect 178567 203869 178601 203897
rect 178629 203869 193899 203897
rect 193927 203869 193961 203897
rect 193989 203869 209259 203897
rect 209287 203869 209321 203897
rect 209349 203869 224619 203897
rect 224647 203869 224681 203897
rect 224709 203869 239979 203897
rect 240007 203869 240041 203897
rect 240069 203869 256437 203897
rect 256465 203869 256499 203897
rect 256527 203869 256561 203897
rect 256589 203869 256623 203897
rect 256651 203869 265437 203897
rect 265465 203869 265499 203897
rect 265527 203869 265561 203897
rect 265589 203869 265623 203897
rect 265651 203869 274437 203897
rect 274465 203869 274499 203897
rect 274527 203869 274561 203897
rect 274589 203869 274623 203897
rect 274651 203869 283437 203897
rect 283465 203869 283499 203897
rect 283527 203869 283561 203897
rect 283589 203869 283623 203897
rect 283651 203869 292437 203897
rect 292465 203869 292499 203897
rect 292527 203869 292561 203897
rect 292589 203869 292623 203897
rect 292651 203869 299736 203897
rect 299764 203869 299798 203897
rect 299826 203869 299860 203897
rect 299888 203869 299922 203897
rect 299950 203869 299998 203897
rect -6 203835 299998 203869
rect -6 203807 42 203835
rect 70 203807 104 203835
rect 132 203807 166 203835
rect 194 203807 228 203835
rect 256 203807 4437 203835
rect 4465 203807 4499 203835
rect 4527 203807 4561 203835
rect 4589 203807 4623 203835
rect 4651 203807 13437 203835
rect 13465 203807 13499 203835
rect 13527 203807 13561 203835
rect 13589 203807 13623 203835
rect 13651 203807 22437 203835
rect 22465 203807 22499 203835
rect 22527 203807 22561 203835
rect 22589 203807 22623 203835
rect 22651 203807 24939 203835
rect 24967 203807 25001 203835
rect 25029 203807 31437 203835
rect 31465 203807 31499 203835
rect 31527 203807 31561 203835
rect 31589 203807 31623 203835
rect 31651 203807 40299 203835
rect 40327 203807 40361 203835
rect 40389 203807 55659 203835
rect 55687 203807 55721 203835
rect 55749 203807 71019 203835
rect 71047 203807 71081 203835
rect 71109 203807 86379 203835
rect 86407 203807 86441 203835
rect 86469 203807 101739 203835
rect 101767 203807 101801 203835
rect 101829 203807 117099 203835
rect 117127 203807 117161 203835
rect 117189 203807 132459 203835
rect 132487 203807 132521 203835
rect 132549 203807 147819 203835
rect 147847 203807 147881 203835
rect 147909 203807 163179 203835
rect 163207 203807 163241 203835
rect 163269 203807 178539 203835
rect 178567 203807 178601 203835
rect 178629 203807 193899 203835
rect 193927 203807 193961 203835
rect 193989 203807 209259 203835
rect 209287 203807 209321 203835
rect 209349 203807 224619 203835
rect 224647 203807 224681 203835
rect 224709 203807 239979 203835
rect 240007 203807 240041 203835
rect 240069 203807 256437 203835
rect 256465 203807 256499 203835
rect 256527 203807 256561 203835
rect 256589 203807 256623 203835
rect 256651 203807 265437 203835
rect 265465 203807 265499 203835
rect 265527 203807 265561 203835
rect 265589 203807 265623 203835
rect 265651 203807 274437 203835
rect 274465 203807 274499 203835
rect 274527 203807 274561 203835
rect 274589 203807 274623 203835
rect 274651 203807 283437 203835
rect 283465 203807 283499 203835
rect 283527 203807 283561 203835
rect 283589 203807 283623 203835
rect 283651 203807 292437 203835
rect 292465 203807 292499 203835
rect 292527 203807 292561 203835
rect 292589 203807 292623 203835
rect 292651 203807 299736 203835
rect 299764 203807 299798 203835
rect 299826 203807 299860 203835
rect 299888 203807 299922 203835
rect 299950 203807 299998 203835
rect -6 203773 299998 203807
rect -6 203745 42 203773
rect 70 203745 104 203773
rect 132 203745 166 203773
rect 194 203745 228 203773
rect 256 203745 4437 203773
rect 4465 203745 4499 203773
rect 4527 203745 4561 203773
rect 4589 203745 4623 203773
rect 4651 203745 13437 203773
rect 13465 203745 13499 203773
rect 13527 203745 13561 203773
rect 13589 203745 13623 203773
rect 13651 203745 22437 203773
rect 22465 203745 22499 203773
rect 22527 203745 22561 203773
rect 22589 203745 22623 203773
rect 22651 203745 24939 203773
rect 24967 203745 25001 203773
rect 25029 203745 31437 203773
rect 31465 203745 31499 203773
rect 31527 203745 31561 203773
rect 31589 203745 31623 203773
rect 31651 203745 40299 203773
rect 40327 203745 40361 203773
rect 40389 203745 55659 203773
rect 55687 203745 55721 203773
rect 55749 203745 71019 203773
rect 71047 203745 71081 203773
rect 71109 203745 86379 203773
rect 86407 203745 86441 203773
rect 86469 203745 101739 203773
rect 101767 203745 101801 203773
rect 101829 203745 117099 203773
rect 117127 203745 117161 203773
rect 117189 203745 132459 203773
rect 132487 203745 132521 203773
rect 132549 203745 147819 203773
rect 147847 203745 147881 203773
rect 147909 203745 163179 203773
rect 163207 203745 163241 203773
rect 163269 203745 178539 203773
rect 178567 203745 178601 203773
rect 178629 203745 193899 203773
rect 193927 203745 193961 203773
rect 193989 203745 209259 203773
rect 209287 203745 209321 203773
rect 209349 203745 224619 203773
rect 224647 203745 224681 203773
rect 224709 203745 239979 203773
rect 240007 203745 240041 203773
rect 240069 203745 256437 203773
rect 256465 203745 256499 203773
rect 256527 203745 256561 203773
rect 256589 203745 256623 203773
rect 256651 203745 265437 203773
rect 265465 203745 265499 203773
rect 265527 203745 265561 203773
rect 265589 203745 265623 203773
rect 265651 203745 274437 203773
rect 274465 203745 274499 203773
rect 274527 203745 274561 203773
rect 274589 203745 274623 203773
rect 274651 203745 283437 203773
rect 283465 203745 283499 203773
rect 283527 203745 283561 203773
rect 283589 203745 283623 203773
rect 283651 203745 292437 203773
rect 292465 203745 292499 203773
rect 292527 203745 292561 203773
rect 292589 203745 292623 203773
rect 292651 203745 299736 203773
rect 299764 203745 299798 203773
rect 299826 203745 299860 203773
rect 299888 203745 299922 203773
rect 299950 203745 299998 203773
rect -6 203697 299998 203745
rect -6 200959 299998 201007
rect -6 200931 522 200959
rect 550 200931 584 200959
rect 612 200931 646 200959
rect 674 200931 708 200959
rect 736 200931 2577 200959
rect 2605 200931 2639 200959
rect 2667 200931 2701 200959
rect 2729 200931 2763 200959
rect 2791 200931 11577 200959
rect 11605 200931 11639 200959
rect 11667 200931 11701 200959
rect 11729 200931 11763 200959
rect 11791 200931 17259 200959
rect 17287 200931 17321 200959
rect 17349 200931 20577 200959
rect 20605 200931 20639 200959
rect 20667 200931 20701 200959
rect 20729 200931 20763 200959
rect 20791 200931 29577 200959
rect 29605 200931 29639 200959
rect 29667 200931 29701 200959
rect 29729 200931 29763 200959
rect 29791 200931 32619 200959
rect 32647 200931 32681 200959
rect 32709 200931 47979 200959
rect 48007 200931 48041 200959
rect 48069 200931 63339 200959
rect 63367 200931 63401 200959
rect 63429 200931 78699 200959
rect 78727 200931 78761 200959
rect 78789 200931 94059 200959
rect 94087 200931 94121 200959
rect 94149 200931 109419 200959
rect 109447 200931 109481 200959
rect 109509 200931 124779 200959
rect 124807 200931 124841 200959
rect 124869 200931 140139 200959
rect 140167 200931 140201 200959
rect 140229 200931 155499 200959
rect 155527 200931 155561 200959
rect 155589 200931 170859 200959
rect 170887 200931 170921 200959
rect 170949 200931 186219 200959
rect 186247 200931 186281 200959
rect 186309 200931 201579 200959
rect 201607 200931 201641 200959
rect 201669 200931 216939 200959
rect 216967 200931 217001 200959
rect 217029 200931 232299 200959
rect 232327 200931 232361 200959
rect 232389 200931 247659 200959
rect 247687 200931 247721 200959
rect 247749 200931 254577 200959
rect 254605 200931 254639 200959
rect 254667 200931 254701 200959
rect 254729 200931 254763 200959
rect 254791 200931 263577 200959
rect 263605 200931 263639 200959
rect 263667 200931 263701 200959
rect 263729 200931 263763 200959
rect 263791 200931 272577 200959
rect 272605 200931 272639 200959
rect 272667 200931 272701 200959
rect 272729 200931 272763 200959
rect 272791 200931 281577 200959
rect 281605 200931 281639 200959
rect 281667 200931 281701 200959
rect 281729 200931 281763 200959
rect 281791 200931 290577 200959
rect 290605 200931 290639 200959
rect 290667 200931 290701 200959
rect 290729 200931 290763 200959
rect 290791 200931 299256 200959
rect 299284 200931 299318 200959
rect 299346 200931 299380 200959
rect 299408 200931 299442 200959
rect 299470 200931 299998 200959
rect -6 200897 299998 200931
rect -6 200869 522 200897
rect 550 200869 584 200897
rect 612 200869 646 200897
rect 674 200869 708 200897
rect 736 200869 2577 200897
rect 2605 200869 2639 200897
rect 2667 200869 2701 200897
rect 2729 200869 2763 200897
rect 2791 200869 11577 200897
rect 11605 200869 11639 200897
rect 11667 200869 11701 200897
rect 11729 200869 11763 200897
rect 11791 200869 17259 200897
rect 17287 200869 17321 200897
rect 17349 200869 20577 200897
rect 20605 200869 20639 200897
rect 20667 200869 20701 200897
rect 20729 200869 20763 200897
rect 20791 200869 29577 200897
rect 29605 200869 29639 200897
rect 29667 200869 29701 200897
rect 29729 200869 29763 200897
rect 29791 200869 32619 200897
rect 32647 200869 32681 200897
rect 32709 200869 47979 200897
rect 48007 200869 48041 200897
rect 48069 200869 63339 200897
rect 63367 200869 63401 200897
rect 63429 200869 78699 200897
rect 78727 200869 78761 200897
rect 78789 200869 94059 200897
rect 94087 200869 94121 200897
rect 94149 200869 109419 200897
rect 109447 200869 109481 200897
rect 109509 200869 124779 200897
rect 124807 200869 124841 200897
rect 124869 200869 140139 200897
rect 140167 200869 140201 200897
rect 140229 200869 155499 200897
rect 155527 200869 155561 200897
rect 155589 200869 170859 200897
rect 170887 200869 170921 200897
rect 170949 200869 186219 200897
rect 186247 200869 186281 200897
rect 186309 200869 201579 200897
rect 201607 200869 201641 200897
rect 201669 200869 216939 200897
rect 216967 200869 217001 200897
rect 217029 200869 232299 200897
rect 232327 200869 232361 200897
rect 232389 200869 247659 200897
rect 247687 200869 247721 200897
rect 247749 200869 254577 200897
rect 254605 200869 254639 200897
rect 254667 200869 254701 200897
rect 254729 200869 254763 200897
rect 254791 200869 263577 200897
rect 263605 200869 263639 200897
rect 263667 200869 263701 200897
rect 263729 200869 263763 200897
rect 263791 200869 272577 200897
rect 272605 200869 272639 200897
rect 272667 200869 272701 200897
rect 272729 200869 272763 200897
rect 272791 200869 281577 200897
rect 281605 200869 281639 200897
rect 281667 200869 281701 200897
rect 281729 200869 281763 200897
rect 281791 200869 290577 200897
rect 290605 200869 290639 200897
rect 290667 200869 290701 200897
rect 290729 200869 290763 200897
rect 290791 200869 299256 200897
rect 299284 200869 299318 200897
rect 299346 200869 299380 200897
rect 299408 200869 299442 200897
rect 299470 200869 299998 200897
rect -6 200835 299998 200869
rect -6 200807 522 200835
rect 550 200807 584 200835
rect 612 200807 646 200835
rect 674 200807 708 200835
rect 736 200807 2577 200835
rect 2605 200807 2639 200835
rect 2667 200807 2701 200835
rect 2729 200807 2763 200835
rect 2791 200807 11577 200835
rect 11605 200807 11639 200835
rect 11667 200807 11701 200835
rect 11729 200807 11763 200835
rect 11791 200807 17259 200835
rect 17287 200807 17321 200835
rect 17349 200807 20577 200835
rect 20605 200807 20639 200835
rect 20667 200807 20701 200835
rect 20729 200807 20763 200835
rect 20791 200807 29577 200835
rect 29605 200807 29639 200835
rect 29667 200807 29701 200835
rect 29729 200807 29763 200835
rect 29791 200807 32619 200835
rect 32647 200807 32681 200835
rect 32709 200807 47979 200835
rect 48007 200807 48041 200835
rect 48069 200807 63339 200835
rect 63367 200807 63401 200835
rect 63429 200807 78699 200835
rect 78727 200807 78761 200835
rect 78789 200807 94059 200835
rect 94087 200807 94121 200835
rect 94149 200807 109419 200835
rect 109447 200807 109481 200835
rect 109509 200807 124779 200835
rect 124807 200807 124841 200835
rect 124869 200807 140139 200835
rect 140167 200807 140201 200835
rect 140229 200807 155499 200835
rect 155527 200807 155561 200835
rect 155589 200807 170859 200835
rect 170887 200807 170921 200835
rect 170949 200807 186219 200835
rect 186247 200807 186281 200835
rect 186309 200807 201579 200835
rect 201607 200807 201641 200835
rect 201669 200807 216939 200835
rect 216967 200807 217001 200835
rect 217029 200807 232299 200835
rect 232327 200807 232361 200835
rect 232389 200807 247659 200835
rect 247687 200807 247721 200835
rect 247749 200807 254577 200835
rect 254605 200807 254639 200835
rect 254667 200807 254701 200835
rect 254729 200807 254763 200835
rect 254791 200807 263577 200835
rect 263605 200807 263639 200835
rect 263667 200807 263701 200835
rect 263729 200807 263763 200835
rect 263791 200807 272577 200835
rect 272605 200807 272639 200835
rect 272667 200807 272701 200835
rect 272729 200807 272763 200835
rect 272791 200807 281577 200835
rect 281605 200807 281639 200835
rect 281667 200807 281701 200835
rect 281729 200807 281763 200835
rect 281791 200807 290577 200835
rect 290605 200807 290639 200835
rect 290667 200807 290701 200835
rect 290729 200807 290763 200835
rect 290791 200807 299256 200835
rect 299284 200807 299318 200835
rect 299346 200807 299380 200835
rect 299408 200807 299442 200835
rect 299470 200807 299998 200835
rect -6 200773 299998 200807
rect -6 200745 522 200773
rect 550 200745 584 200773
rect 612 200745 646 200773
rect 674 200745 708 200773
rect 736 200745 2577 200773
rect 2605 200745 2639 200773
rect 2667 200745 2701 200773
rect 2729 200745 2763 200773
rect 2791 200745 11577 200773
rect 11605 200745 11639 200773
rect 11667 200745 11701 200773
rect 11729 200745 11763 200773
rect 11791 200745 17259 200773
rect 17287 200745 17321 200773
rect 17349 200745 20577 200773
rect 20605 200745 20639 200773
rect 20667 200745 20701 200773
rect 20729 200745 20763 200773
rect 20791 200745 29577 200773
rect 29605 200745 29639 200773
rect 29667 200745 29701 200773
rect 29729 200745 29763 200773
rect 29791 200745 32619 200773
rect 32647 200745 32681 200773
rect 32709 200745 47979 200773
rect 48007 200745 48041 200773
rect 48069 200745 63339 200773
rect 63367 200745 63401 200773
rect 63429 200745 78699 200773
rect 78727 200745 78761 200773
rect 78789 200745 94059 200773
rect 94087 200745 94121 200773
rect 94149 200745 109419 200773
rect 109447 200745 109481 200773
rect 109509 200745 124779 200773
rect 124807 200745 124841 200773
rect 124869 200745 140139 200773
rect 140167 200745 140201 200773
rect 140229 200745 155499 200773
rect 155527 200745 155561 200773
rect 155589 200745 170859 200773
rect 170887 200745 170921 200773
rect 170949 200745 186219 200773
rect 186247 200745 186281 200773
rect 186309 200745 201579 200773
rect 201607 200745 201641 200773
rect 201669 200745 216939 200773
rect 216967 200745 217001 200773
rect 217029 200745 232299 200773
rect 232327 200745 232361 200773
rect 232389 200745 247659 200773
rect 247687 200745 247721 200773
rect 247749 200745 254577 200773
rect 254605 200745 254639 200773
rect 254667 200745 254701 200773
rect 254729 200745 254763 200773
rect 254791 200745 263577 200773
rect 263605 200745 263639 200773
rect 263667 200745 263701 200773
rect 263729 200745 263763 200773
rect 263791 200745 272577 200773
rect 272605 200745 272639 200773
rect 272667 200745 272701 200773
rect 272729 200745 272763 200773
rect 272791 200745 281577 200773
rect 281605 200745 281639 200773
rect 281667 200745 281701 200773
rect 281729 200745 281763 200773
rect 281791 200745 290577 200773
rect 290605 200745 290639 200773
rect 290667 200745 290701 200773
rect 290729 200745 290763 200773
rect 290791 200745 299256 200773
rect 299284 200745 299318 200773
rect 299346 200745 299380 200773
rect 299408 200745 299442 200773
rect 299470 200745 299998 200773
rect -6 200697 299998 200745
rect -6 194959 299998 195007
rect -6 194931 42 194959
rect 70 194931 104 194959
rect 132 194931 166 194959
rect 194 194931 228 194959
rect 256 194931 4437 194959
rect 4465 194931 4499 194959
rect 4527 194931 4561 194959
rect 4589 194931 4623 194959
rect 4651 194931 13437 194959
rect 13465 194931 13499 194959
rect 13527 194931 13561 194959
rect 13589 194931 13623 194959
rect 13651 194931 22437 194959
rect 22465 194931 22499 194959
rect 22527 194931 22561 194959
rect 22589 194931 22623 194959
rect 22651 194931 24939 194959
rect 24967 194931 25001 194959
rect 25029 194931 31437 194959
rect 31465 194931 31499 194959
rect 31527 194931 31561 194959
rect 31589 194931 31623 194959
rect 31651 194931 40299 194959
rect 40327 194931 40361 194959
rect 40389 194931 55659 194959
rect 55687 194931 55721 194959
rect 55749 194931 71019 194959
rect 71047 194931 71081 194959
rect 71109 194931 86379 194959
rect 86407 194931 86441 194959
rect 86469 194931 101739 194959
rect 101767 194931 101801 194959
rect 101829 194931 117099 194959
rect 117127 194931 117161 194959
rect 117189 194931 132459 194959
rect 132487 194931 132521 194959
rect 132549 194931 147819 194959
rect 147847 194931 147881 194959
rect 147909 194931 163179 194959
rect 163207 194931 163241 194959
rect 163269 194931 178539 194959
rect 178567 194931 178601 194959
rect 178629 194931 193899 194959
rect 193927 194931 193961 194959
rect 193989 194931 209259 194959
rect 209287 194931 209321 194959
rect 209349 194931 224619 194959
rect 224647 194931 224681 194959
rect 224709 194931 239979 194959
rect 240007 194931 240041 194959
rect 240069 194931 256437 194959
rect 256465 194931 256499 194959
rect 256527 194931 256561 194959
rect 256589 194931 256623 194959
rect 256651 194931 265437 194959
rect 265465 194931 265499 194959
rect 265527 194931 265561 194959
rect 265589 194931 265623 194959
rect 265651 194931 274437 194959
rect 274465 194931 274499 194959
rect 274527 194931 274561 194959
rect 274589 194931 274623 194959
rect 274651 194931 283437 194959
rect 283465 194931 283499 194959
rect 283527 194931 283561 194959
rect 283589 194931 283623 194959
rect 283651 194931 292437 194959
rect 292465 194931 292499 194959
rect 292527 194931 292561 194959
rect 292589 194931 292623 194959
rect 292651 194931 299736 194959
rect 299764 194931 299798 194959
rect 299826 194931 299860 194959
rect 299888 194931 299922 194959
rect 299950 194931 299998 194959
rect -6 194897 299998 194931
rect -6 194869 42 194897
rect 70 194869 104 194897
rect 132 194869 166 194897
rect 194 194869 228 194897
rect 256 194869 4437 194897
rect 4465 194869 4499 194897
rect 4527 194869 4561 194897
rect 4589 194869 4623 194897
rect 4651 194869 13437 194897
rect 13465 194869 13499 194897
rect 13527 194869 13561 194897
rect 13589 194869 13623 194897
rect 13651 194869 22437 194897
rect 22465 194869 22499 194897
rect 22527 194869 22561 194897
rect 22589 194869 22623 194897
rect 22651 194869 24939 194897
rect 24967 194869 25001 194897
rect 25029 194869 31437 194897
rect 31465 194869 31499 194897
rect 31527 194869 31561 194897
rect 31589 194869 31623 194897
rect 31651 194869 40299 194897
rect 40327 194869 40361 194897
rect 40389 194869 55659 194897
rect 55687 194869 55721 194897
rect 55749 194869 71019 194897
rect 71047 194869 71081 194897
rect 71109 194869 86379 194897
rect 86407 194869 86441 194897
rect 86469 194869 101739 194897
rect 101767 194869 101801 194897
rect 101829 194869 117099 194897
rect 117127 194869 117161 194897
rect 117189 194869 132459 194897
rect 132487 194869 132521 194897
rect 132549 194869 147819 194897
rect 147847 194869 147881 194897
rect 147909 194869 163179 194897
rect 163207 194869 163241 194897
rect 163269 194869 178539 194897
rect 178567 194869 178601 194897
rect 178629 194869 193899 194897
rect 193927 194869 193961 194897
rect 193989 194869 209259 194897
rect 209287 194869 209321 194897
rect 209349 194869 224619 194897
rect 224647 194869 224681 194897
rect 224709 194869 239979 194897
rect 240007 194869 240041 194897
rect 240069 194869 256437 194897
rect 256465 194869 256499 194897
rect 256527 194869 256561 194897
rect 256589 194869 256623 194897
rect 256651 194869 265437 194897
rect 265465 194869 265499 194897
rect 265527 194869 265561 194897
rect 265589 194869 265623 194897
rect 265651 194869 274437 194897
rect 274465 194869 274499 194897
rect 274527 194869 274561 194897
rect 274589 194869 274623 194897
rect 274651 194869 283437 194897
rect 283465 194869 283499 194897
rect 283527 194869 283561 194897
rect 283589 194869 283623 194897
rect 283651 194869 292437 194897
rect 292465 194869 292499 194897
rect 292527 194869 292561 194897
rect 292589 194869 292623 194897
rect 292651 194869 299736 194897
rect 299764 194869 299798 194897
rect 299826 194869 299860 194897
rect 299888 194869 299922 194897
rect 299950 194869 299998 194897
rect -6 194835 299998 194869
rect -6 194807 42 194835
rect 70 194807 104 194835
rect 132 194807 166 194835
rect 194 194807 228 194835
rect 256 194807 4437 194835
rect 4465 194807 4499 194835
rect 4527 194807 4561 194835
rect 4589 194807 4623 194835
rect 4651 194807 13437 194835
rect 13465 194807 13499 194835
rect 13527 194807 13561 194835
rect 13589 194807 13623 194835
rect 13651 194807 22437 194835
rect 22465 194807 22499 194835
rect 22527 194807 22561 194835
rect 22589 194807 22623 194835
rect 22651 194807 24939 194835
rect 24967 194807 25001 194835
rect 25029 194807 31437 194835
rect 31465 194807 31499 194835
rect 31527 194807 31561 194835
rect 31589 194807 31623 194835
rect 31651 194807 40299 194835
rect 40327 194807 40361 194835
rect 40389 194807 55659 194835
rect 55687 194807 55721 194835
rect 55749 194807 71019 194835
rect 71047 194807 71081 194835
rect 71109 194807 86379 194835
rect 86407 194807 86441 194835
rect 86469 194807 101739 194835
rect 101767 194807 101801 194835
rect 101829 194807 117099 194835
rect 117127 194807 117161 194835
rect 117189 194807 132459 194835
rect 132487 194807 132521 194835
rect 132549 194807 147819 194835
rect 147847 194807 147881 194835
rect 147909 194807 163179 194835
rect 163207 194807 163241 194835
rect 163269 194807 178539 194835
rect 178567 194807 178601 194835
rect 178629 194807 193899 194835
rect 193927 194807 193961 194835
rect 193989 194807 209259 194835
rect 209287 194807 209321 194835
rect 209349 194807 224619 194835
rect 224647 194807 224681 194835
rect 224709 194807 239979 194835
rect 240007 194807 240041 194835
rect 240069 194807 256437 194835
rect 256465 194807 256499 194835
rect 256527 194807 256561 194835
rect 256589 194807 256623 194835
rect 256651 194807 265437 194835
rect 265465 194807 265499 194835
rect 265527 194807 265561 194835
rect 265589 194807 265623 194835
rect 265651 194807 274437 194835
rect 274465 194807 274499 194835
rect 274527 194807 274561 194835
rect 274589 194807 274623 194835
rect 274651 194807 283437 194835
rect 283465 194807 283499 194835
rect 283527 194807 283561 194835
rect 283589 194807 283623 194835
rect 283651 194807 292437 194835
rect 292465 194807 292499 194835
rect 292527 194807 292561 194835
rect 292589 194807 292623 194835
rect 292651 194807 299736 194835
rect 299764 194807 299798 194835
rect 299826 194807 299860 194835
rect 299888 194807 299922 194835
rect 299950 194807 299998 194835
rect -6 194773 299998 194807
rect -6 194745 42 194773
rect 70 194745 104 194773
rect 132 194745 166 194773
rect 194 194745 228 194773
rect 256 194745 4437 194773
rect 4465 194745 4499 194773
rect 4527 194745 4561 194773
rect 4589 194745 4623 194773
rect 4651 194745 13437 194773
rect 13465 194745 13499 194773
rect 13527 194745 13561 194773
rect 13589 194745 13623 194773
rect 13651 194745 22437 194773
rect 22465 194745 22499 194773
rect 22527 194745 22561 194773
rect 22589 194745 22623 194773
rect 22651 194745 24939 194773
rect 24967 194745 25001 194773
rect 25029 194745 31437 194773
rect 31465 194745 31499 194773
rect 31527 194745 31561 194773
rect 31589 194745 31623 194773
rect 31651 194745 40299 194773
rect 40327 194745 40361 194773
rect 40389 194745 55659 194773
rect 55687 194745 55721 194773
rect 55749 194745 71019 194773
rect 71047 194745 71081 194773
rect 71109 194745 86379 194773
rect 86407 194745 86441 194773
rect 86469 194745 101739 194773
rect 101767 194745 101801 194773
rect 101829 194745 117099 194773
rect 117127 194745 117161 194773
rect 117189 194745 132459 194773
rect 132487 194745 132521 194773
rect 132549 194745 147819 194773
rect 147847 194745 147881 194773
rect 147909 194745 163179 194773
rect 163207 194745 163241 194773
rect 163269 194745 178539 194773
rect 178567 194745 178601 194773
rect 178629 194745 193899 194773
rect 193927 194745 193961 194773
rect 193989 194745 209259 194773
rect 209287 194745 209321 194773
rect 209349 194745 224619 194773
rect 224647 194745 224681 194773
rect 224709 194745 239979 194773
rect 240007 194745 240041 194773
rect 240069 194745 256437 194773
rect 256465 194745 256499 194773
rect 256527 194745 256561 194773
rect 256589 194745 256623 194773
rect 256651 194745 265437 194773
rect 265465 194745 265499 194773
rect 265527 194745 265561 194773
rect 265589 194745 265623 194773
rect 265651 194745 274437 194773
rect 274465 194745 274499 194773
rect 274527 194745 274561 194773
rect 274589 194745 274623 194773
rect 274651 194745 283437 194773
rect 283465 194745 283499 194773
rect 283527 194745 283561 194773
rect 283589 194745 283623 194773
rect 283651 194745 292437 194773
rect 292465 194745 292499 194773
rect 292527 194745 292561 194773
rect 292589 194745 292623 194773
rect 292651 194745 299736 194773
rect 299764 194745 299798 194773
rect 299826 194745 299860 194773
rect 299888 194745 299922 194773
rect 299950 194745 299998 194773
rect -6 194697 299998 194745
rect -6 191959 299998 192007
rect -6 191931 522 191959
rect 550 191931 584 191959
rect 612 191931 646 191959
rect 674 191931 708 191959
rect 736 191931 2577 191959
rect 2605 191931 2639 191959
rect 2667 191931 2701 191959
rect 2729 191931 2763 191959
rect 2791 191931 11577 191959
rect 11605 191931 11639 191959
rect 11667 191931 11701 191959
rect 11729 191931 11763 191959
rect 11791 191931 17259 191959
rect 17287 191931 17321 191959
rect 17349 191931 20577 191959
rect 20605 191931 20639 191959
rect 20667 191931 20701 191959
rect 20729 191931 20763 191959
rect 20791 191931 29577 191959
rect 29605 191931 29639 191959
rect 29667 191931 29701 191959
rect 29729 191931 29763 191959
rect 29791 191931 32619 191959
rect 32647 191931 32681 191959
rect 32709 191931 47979 191959
rect 48007 191931 48041 191959
rect 48069 191931 63339 191959
rect 63367 191931 63401 191959
rect 63429 191931 78699 191959
rect 78727 191931 78761 191959
rect 78789 191931 94059 191959
rect 94087 191931 94121 191959
rect 94149 191931 109419 191959
rect 109447 191931 109481 191959
rect 109509 191931 124779 191959
rect 124807 191931 124841 191959
rect 124869 191931 140139 191959
rect 140167 191931 140201 191959
rect 140229 191931 155499 191959
rect 155527 191931 155561 191959
rect 155589 191931 170859 191959
rect 170887 191931 170921 191959
rect 170949 191931 186219 191959
rect 186247 191931 186281 191959
rect 186309 191931 201579 191959
rect 201607 191931 201641 191959
rect 201669 191931 216939 191959
rect 216967 191931 217001 191959
rect 217029 191931 232299 191959
rect 232327 191931 232361 191959
rect 232389 191931 247659 191959
rect 247687 191931 247721 191959
rect 247749 191931 254577 191959
rect 254605 191931 254639 191959
rect 254667 191931 254701 191959
rect 254729 191931 254763 191959
rect 254791 191931 263577 191959
rect 263605 191931 263639 191959
rect 263667 191931 263701 191959
rect 263729 191931 263763 191959
rect 263791 191931 272577 191959
rect 272605 191931 272639 191959
rect 272667 191931 272701 191959
rect 272729 191931 272763 191959
rect 272791 191931 281577 191959
rect 281605 191931 281639 191959
rect 281667 191931 281701 191959
rect 281729 191931 281763 191959
rect 281791 191931 290577 191959
rect 290605 191931 290639 191959
rect 290667 191931 290701 191959
rect 290729 191931 290763 191959
rect 290791 191931 299256 191959
rect 299284 191931 299318 191959
rect 299346 191931 299380 191959
rect 299408 191931 299442 191959
rect 299470 191931 299998 191959
rect -6 191897 299998 191931
rect -6 191869 522 191897
rect 550 191869 584 191897
rect 612 191869 646 191897
rect 674 191869 708 191897
rect 736 191869 2577 191897
rect 2605 191869 2639 191897
rect 2667 191869 2701 191897
rect 2729 191869 2763 191897
rect 2791 191869 11577 191897
rect 11605 191869 11639 191897
rect 11667 191869 11701 191897
rect 11729 191869 11763 191897
rect 11791 191869 17259 191897
rect 17287 191869 17321 191897
rect 17349 191869 20577 191897
rect 20605 191869 20639 191897
rect 20667 191869 20701 191897
rect 20729 191869 20763 191897
rect 20791 191869 29577 191897
rect 29605 191869 29639 191897
rect 29667 191869 29701 191897
rect 29729 191869 29763 191897
rect 29791 191869 32619 191897
rect 32647 191869 32681 191897
rect 32709 191869 47979 191897
rect 48007 191869 48041 191897
rect 48069 191869 63339 191897
rect 63367 191869 63401 191897
rect 63429 191869 78699 191897
rect 78727 191869 78761 191897
rect 78789 191869 94059 191897
rect 94087 191869 94121 191897
rect 94149 191869 109419 191897
rect 109447 191869 109481 191897
rect 109509 191869 124779 191897
rect 124807 191869 124841 191897
rect 124869 191869 140139 191897
rect 140167 191869 140201 191897
rect 140229 191869 155499 191897
rect 155527 191869 155561 191897
rect 155589 191869 170859 191897
rect 170887 191869 170921 191897
rect 170949 191869 186219 191897
rect 186247 191869 186281 191897
rect 186309 191869 201579 191897
rect 201607 191869 201641 191897
rect 201669 191869 216939 191897
rect 216967 191869 217001 191897
rect 217029 191869 232299 191897
rect 232327 191869 232361 191897
rect 232389 191869 247659 191897
rect 247687 191869 247721 191897
rect 247749 191869 254577 191897
rect 254605 191869 254639 191897
rect 254667 191869 254701 191897
rect 254729 191869 254763 191897
rect 254791 191869 263577 191897
rect 263605 191869 263639 191897
rect 263667 191869 263701 191897
rect 263729 191869 263763 191897
rect 263791 191869 272577 191897
rect 272605 191869 272639 191897
rect 272667 191869 272701 191897
rect 272729 191869 272763 191897
rect 272791 191869 281577 191897
rect 281605 191869 281639 191897
rect 281667 191869 281701 191897
rect 281729 191869 281763 191897
rect 281791 191869 290577 191897
rect 290605 191869 290639 191897
rect 290667 191869 290701 191897
rect 290729 191869 290763 191897
rect 290791 191869 299256 191897
rect 299284 191869 299318 191897
rect 299346 191869 299380 191897
rect 299408 191869 299442 191897
rect 299470 191869 299998 191897
rect -6 191835 299998 191869
rect -6 191807 522 191835
rect 550 191807 584 191835
rect 612 191807 646 191835
rect 674 191807 708 191835
rect 736 191807 2577 191835
rect 2605 191807 2639 191835
rect 2667 191807 2701 191835
rect 2729 191807 2763 191835
rect 2791 191807 11577 191835
rect 11605 191807 11639 191835
rect 11667 191807 11701 191835
rect 11729 191807 11763 191835
rect 11791 191807 17259 191835
rect 17287 191807 17321 191835
rect 17349 191807 20577 191835
rect 20605 191807 20639 191835
rect 20667 191807 20701 191835
rect 20729 191807 20763 191835
rect 20791 191807 29577 191835
rect 29605 191807 29639 191835
rect 29667 191807 29701 191835
rect 29729 191807 29763 191835
rect 29791 191807 32619 191835
rect 32647 191807 32681 191835
rect 32709 191807 47979 191835
rect 48007 191807 48041 191835
rect 48069 191807 63339 191835
rect 63367 191807 63401 191835
rect 63429 191807 78699 191835
rect 78727 191807 78761 191835
rect 78789 191807 94059 191835
rect 94087 191807 94121 191835
rect 94149 191807 109419 191835
rect 109447 191807 109481 191835
rect 109509 191807 124779 191835
rect 124807 191807 124841 191835
rect 124869 191807 140139 191835
rect 140167 191807 140201 191835
rect 140229 191807 155499 191835
rect 155527 191807 155561 191835
rect 155589 191807 170859 191835
rect 170887 191807 170921 191835
rect 170949 191807 186219 191835
rect 186247 191807 186281 191835
rect 186309 191807 201579 191835
rect 201607 191807 201641 191835
rect 201669 191807 216939 191835
rect 216967 191807 217001 191835
rect 217029 191807 232299 191835
rect 232327 191807 232361 191835
rect 232389 191807 247659 191835
rect 247687 191807 247721 191835
rect 247749 191807 254577 191835
rect 254605 191807 254639 191835
rect 254667 191807 254701 191835
rect 254729 191807 254763 191835
rect 254791 191807 263577 191835
rect 263605 191807 263639 191835
rect 263667 191807 263701 191835
rect 263729 191807 263763 191835
rect 263791 191807 272577 191835
rect 272605 191807 272639 191835
rect 272667 191807 272701 191835
rect 272729 191807 272763 191835
rect 272791 191807 281577 191835
rect 281605 191807 281639 191835
rect 281667 191807 281701 191835
rect 281729 191807 281763 191835
rect 281791 191807 290577 191835
rect 290605 191807 290639 191835
rect 290667 191807 290701 191835
rect 290729 191807 290763 191835
rect 290791 191807 299256 191835
rect 299284 191807 299318 191835
rect 299346 191807 299380 191835
rect 299408 191807 299442 191835
rect 299470 191807 299998 191835
rect -6 191773 299998 191807
rect -6 191745 522 191773
rect 550 191745 584 191773
rect 612 191745 646 191773
rect 674 191745 708 191773
rect 736 191745 2577 191773
rect 2605 191745 2639 191773
rect 2667 191745 2701 191773
rect 2729 191745 2763 191773
rect 2791 191745 11577 191773
rect 11605 191745 11639 191773
rect 11667 191745 11701 191773
rect 11729 191745 11763 191773
rect 11791 191745 17259 191773
rect 17287 191745 17321 191773
rect 17349 191745 20577 191773
rect 20605 191745 20639 191773
rect 20667 191745 20701 191773
rect 20729 191745 20763 191773
rect 20791 191745 29577 191773
rect 29605 191745 29639 191773
rect 29667 191745 29701 191773
rect 29729 191745 29763 191773
rect 29791 191745 32619 191773
rect 32647 191745 32681 191773
rect 32709 191745 47979 191773
rect 48007 191745 48041 191773
rect 48069 191745 63339 191773
rect 63367 191745 63401 191773
rect 63429 191745 78699 191773
rect 78727 191745 78761 191773
rect 78789 191745 94059 191773
rect 94087 191745 94121 191773
rect 94149 191745 109419 191773
rect 109447 191745 109481 191773
rect 109509 191745 124779 191773
rect 124807 191745 124841 191773
rect 124869 191745 140139 191773
rect 140167 191745 140201 191773
rect 140229 191745 155499 191773
rect 155527 191745 155561 191773
rect 155589 191745 170859 191773
rect 170887 191745 170921 191773
rect 170949 191745 186219 191773
rect 186247 191745 186281 191773
rect 186309 191745 201579 191773
rect 201607 191745 201641 191773
rect 201669 191745 216939 191773
rect 216967 191745 217001 191773
rect 217029 191745 232299 191773
rect 232327 191745 232361 191773
rect 232389 191745 247659 191773
rect 247687 191745 247721 191773
rect 247749 191745 254577 191773
rect 254605 191745 254639 191773
rect 254667 191745 254701 191773
rect 254729 191745 254763 191773
rect 254791 191745 263577 191773
rect 263605 191745 263639 191773
rect 263667 191745 263701 191773
rect 263729 191745 263763 191773
rect 263791 191745 272577 191773
rect 272605 191745 272639 191773
rect 272667 191745 272701 191773
rect 272729 191745 272763 191773
rect 272791 191745 281577 191773
rect 281605 191745 281639 191773
rect 281667 191745 281701 191773
rect 281729 191745 281763 191773
rect 281791 191745 290577 191773
rect 290605 191745 290639 191773
rect 290667 191745 290701 191773
rect 290729 191745 290763 191773
rect 290791 191745 299256 191773
rect 299284 191745 299318 191773
rect 299346 191745 299380 191773
rect 299408 191745 299442 191773
rect 299470 191745 299998 191773
rect -6 191697 299998 191745
rect -6 185959 299998 186007
rect -6 185931 42 185959
rect 70 185931 104 185959
rect 132 185931 166 185959
rect 194 185931 228 185959
rect 256 185931 4437 185959
rect 4465 185931 4499 185959
rect 4527 185931 4561 185959
rect 4589 185931 4623 185959
rect 4651 185931 13437 185959
rect 13465 185931 13499 185959
rect 13527 185931 13561 185959
rect 13589 185931 13623 185959
rect 13651 185931 22437 185959
rect 22465 185931 22499 185959
rect 22527 185931 22561 185959
rect 22589 185931 22623 185959
rect 22651 185931 24939 185959
rect 24967 185931 25001 185959
rect 25029 185931 31437 185959
rect 31465 185931 31499 185959
rect 31527 185931 31561 185959
rect 31589 185931 31623 185959
rect 31651 185931 40299 185959
rect 40327 185931 40361 185959
rect 40389 185931 55659 185959
rect 55687 185931 55721 185959
rect 55749 185931 71019 185959
rect 71047 185931 71081 185959
rect 71109 185931 86379 185959
rect 86407 185931 86441 185959
rect 86469 185931 101739 185959
rect 101767 185931 101801 185959
rect 101829 185931 117099 185959
rect 117127 185931 117161 185959
rect 117189 185931 132459 185959
rect 132487 185931 132521 185959
rect 132549 185931 147819 185959
rect 147847 185931 147881 185959
rect 147909 185931 163179 185959
rect 163207 185931 163241 185959
rect 163269 185931 178539 185959
rect 178567 185931 178601 185959
rect 178629 185931 193899 185959
rect 193927 185931 193961 185959
rect 193989 185931 209259 185959
rect 209287 185931 209321 185959
rect 209349 185931 224619 185959
rect 224647 185931 224681 185959
rect 224709 185931 239979 185959
rect 240007 185931 240041 185959
rect 240069 185931 256437 185959
rect 256465 185931 256499 185959
rect 256527 185931 256561 185959
rect 256589 185931 256623 185959
rect 256651 185931 265437 185959
rect 265465 185931 265499 185959
rect 265527 185931 265561 185959
rect 265589 185931 265623 185959
rect 265651 185931 274437 185959
rect 274465 185931 274499 185959
rect 274527 185931 274561 185959
rect 274589 185931 274623 185959
rect 274651 185931 283437 185959
rect 283465 185931 283499 185959
rect 283527 185931 283561 185959
rect 283589 185931 283623 185959
rect 283651 185931 292437 185959
rect 292465 185931 292499 185959
rect 292527 185931 292561 185959
rect 292589 185931 292623 185959
rect 292651 185931 299736 185959
rect 299764 185931 299798 185959
rect 299826 185931 299860 185959
rect 299888 185931 299922 185959
rect 299950 185931 299998 185959
rect -6 185897 299998 185931
rect -6 185869 42 185897
rect 70 185869 104 185897
rect 132 185869 166 185897
rect 194 185869 228 185897
rect 256 185869 4437 185897
rect 4465 185869 4499 185897
rect 4527 185869 4561 185897
rect 4589 185869 4623 185897
rect 4651 185869 13437 185897
rect 13465 185869 13499 185897
rect 13527 185869 13561 185897
rect 13589 185869 13623 185897
rect 13651 185869 22437 185897
rect 22465 185869 22499 185897
rect 22527 185869 22561 185897
rect 22589 185869 22623 185897
rect 22651 185869 24939 185897
rect 24967 185869 25001 185897
rect 25029 185869 31437 185897
rect 31465 185869 31499 185897
rect 31527 185869 31561 185897
rect 31589 185869 31623 185897
rect 31651 185869 40299 185897
rect 40327 185869 40361 185897
rect 40389 185869 55659 185897
rect 55687 185869 55721 185897
rect 55749 185869 71019 185897
rect 71047 185869 71081 185897
rect 71109 185869 86379 185897
rect 86407 185869 86441 185897
rect 86469 185869 101739 185897
rect 101767 185869 101801 185897
rect 101829 185869 117099 185897
rect 117127 185869 117161 185897
rect 117189 185869 132459 185897
rect 132487 185869 132521 185897
rect 132549 185869 147819 185897
rect 147847 185869 147881 185897
rect 147909 185869 163179 185897
rect 163207 185869 163241 185897
rect 163269 185869 178539 185897
rect 178567 185869 178601 185897
rect 178629 185869 193899 185897
rect 193927 185869 193961 185897
rect 193989 185869 209259 185897
rect 209287 185869 209321 185897
rect 209349 185869 224619 185897
rect 224647 185869 224681 185897
rect 224709 185869 239979 185897
rect 240007 185869 240041 185897
rect 240069 185869 256437 185897
rect 256465 185869 256499 185897
rect 256527 185869 256561 185897
rect 256589 185869 256623 185897
rect 256651 185869 265437 185897
rect 265465 185869 265499 185897
rect 265527 185869 265561 185897
rect 265589 185869 265623 185897
rect 265651 185869 274437 185897
rect 274465 185869 274499 185897
rect 274527 185869 274561 185897
rect 274589 185869 274623 185897
rect 274651 185869 283437 185897
rect 283465 185869 283499 185897
rect 283527 185869 283561 185897
rect 283589 185869 283623 185897
rect 283651 185869 292437 185897
rect 292465 185869 292499 185897
rect 292527 185869 292561 185897
rect 292589 185869 292623 185897
rect 292651 185869 299736 185897
rect 299764 185869 299798 185897
rect 299826 185869 299860 185897
rect 299888 185869 299922 185897
rect 299950 185869 299998 185897
rect -6 185835 299998 185869
rect -6 185807 42 185835
rect 70 185807 104 185835
rect 132 185807 166 185835
rect 194 185807 228 185835
rect 256 185807 4437 185835
rect 4465 185807 4499 185835
rect 4527 185807 4561 185835
rect 4589 185807 4623 185835
rect 4651 185807 13437 185835
rect 13465 185807 13499 185835
rect 13527 185807 13561 185835
rect 13589 185807 13623 185835
rect 13651 185807 22437 185835
rect 22465 185807 22499 185835
rect 22527 185807 22561 185835
rect 22589 185807 22623 185835
rect 22651 185807 24939 185835
rect 24967 185807 25001 185835
rect 25029 185807 31437 185835
rect 31465 185807 31499 185835
rect 31527 185807 31561 185835
rect 31589 185807 31623 185835
rect 31651 185807 40299 185835
rect 40327 185807 40361 185835
rect 40389 185807 55659 185835
rect 55687 185807 55721 185835
rect 55749 185807 71019 185835
rect 71047 185807 71081 185835
rect 71109 185807 86379 185835
rect 86407 185807 86441 185835
rect 86469 185807 101739 185835
rect 101767 185807 101801 185835
rect 101829 185807 117099 185835
rect 117127 185807 117161 185835
rect 117189 185807 132459 185835
rect 132487 185807 132521 185835
rect 132549 185807 147819 185835
rect 147847 185807 147881 185835
rect 147909 185807 163179 185835
rect 163207 185807 163241 185835
rect 163269 185807 178539 185835
rect 178567 185807 178601 185835
rect 178629 185807 193899 185835
rect 193927 185807 193961 185835
rect 193989 185807 209259 185835
rect 209287 185807 209321 185835
rect 209349 185807 224619 185835
rect 224647 185807 224681 185835
rect 224709 185807 239979 185835
rect 240007 185807 240041 185835
rect 240069 185807 256437 185835
rect 256465 185807 256499 185835
rect 256527 185807 256561 185835
rect 256589 185807 256623 185835
rect 256651 185807 265437 185835
rect 265465 185807 265499 185835
rect 265527 185807 265561 185835
rect 265589 185807 265623 185835
rect 265651 185807 274437 185835
rect 274465 185807 274499 185835
rect 274527 185807 274561 185835
rect 274589 185807 274623 185835
rect 274651 185807 283437 185835
rect 283465 185807 283499 185835
rect 283527 185807 283561 185835
rect 283589 185807 283623 185835
rect 283651 185807 292437 185835
rect 292465 185807 292499 185835
rect 292527 185807 292561 185835
rect 292589 185807 292623 185835
rect 292651 185807 299736 185835
rect 299764 185807 299798 185835
rect 299826 185807 299860 185835
rect 299888 185807 299922 185835
rect 299950 185807 299998 185835
rect -6 185773 299998 185807
rect -6 185745 42 185773
rect 70 185745 104 185773
rect 132 185745 166 185773
rect 194 185745 228 185773
rect 256 185745 4437 185773
rect 4465 185745 4499 185773
rect 4527 185745 4561 185773
rect 4589 185745 4623 185773
rect 4651 185745 13437 185773
rect 13465 185745 13499 185773
rect 13527 185745 13561 185773
rect 13589 185745 13623 185773
rect 13651 185745 22437 185773
rect 22465 185745 22499 185773
rect 22527 185745 22561 185773
rect 22589 185745 22623 185773
rect 22651 185745 24939 185773
rect 24967 185745 25001 185773
rect 25029 185745 31437 185773
rect 31465 185745 31499 185773
rect 31527 185745 31561 185773
rect 31589 185745 31623 185773
rect 31651 185745 40299 185773
rect 40327 185745 40361 185773
rect 40389 185745 55659 185773
rect 55687 185745 55721 185773
rect 55749 185745 71019 185773
rect 71047 185745 71081 185773
rect 71109 185745 86379 185773
rect 86407 185745 86441 185773
rect 86469 185745 101739 185773
rect 101767 185745 101801 185773
rect 101829 185745 117099 185773
rect 117127 185745 117161 185773
rect 117189 185745 132459 185773
rect 132487 185745 132521 185773
rect 132549 185745 147819 185773
rect 147847 185745 147881 185773
rect 147909 185745 163179 185773
rect 163207 185745 163241 185773
rect 163269 185745 178539 185773
rect 178567 185745 178601 185773
rect 178629 185745 193899 185773
rect 193927 185745 193961 185773
rect 193989 185745 209259 185773
rect 209287 185745 209321 185773
rect 209349 185745 224619 185773
rect 224647 185745 224681 185773
rect 224709 185745 239979 185773
rect 240007 185745 240041 185773
rect 240069 185745 256437 185773
rect 256465 185745 256499 185773
rect 256527 185745 256561 185773
rect 256589 185745 256623 185773
rect 256651 185745 265437 185773
rect 265465 185745 265499 185773
rect 265527 185745 265561 185773
rect 265589 185745 265623 185773
rect 265651 185745 274437 185773
rect 274465 185745 274499 185773
rect 274527 185745 274561 185773
rect 274589 185745 274623 185773
rect 274651 185745 283437 185773
rect 283465 185745 283499 185773
rect 283527 185745 283561 185773
rect 283589 185745 283623 185773
rect 283651 185745 292437 185773
rect 292465 185745 292499 185773
rect 292527 185745 292561 185773
rect 292589 185745 292623 185773
rect 292651 185745 299736 185773
rect 299764 185745 299798 185773
rect 299826 185745 299860 185773
rect 299888 185745 299922 185773
rect 299950 185745 299998 185773
rect -6 185697 299998 185745
rect -6 182959 299998 183007
rect -6 182931 522 182959
rect 550 182931 584 182959
rect 612 182931 646 182959
rect 674 182931 708 182959
rect 736 182931 2577 182959
rect 2605 182931 2639 182959
rect 2667 182931 2701 182959
rect 2729 182931 2763 182959
rect 2791 182931 11577 182959
rect 11605 182931 11639 182959
rect 11667 182931 11701 182959
rect 11729 182931 11763 182959
rect 11791 182931 17259 182959
rect 17287 182931 17321 182959
rect 17349 182931 20577 182959
rect 20605 182931 20639 182959
rect 20667 182931 20701 182959
rect 20729 182931 20763 182959
rect 20791 182931 29577 182959
rect 29605 182931 29639 182959
rect 29667 182931 29701 182959
rect 29729 182931 29763 182959
rect 29791 182931 32619 182959
rect 32647 182931 32681 182959
rect 32709 182931 47979 182959
rect 48007 182931 48041 182959
rect 48069 182931 63339 182959
rect 63367 182931 63401 182959
rect 63429 182931 78699 182959
rect 78727 182931 78761 182959
rect 78789 182931 94059 182959
rect 94087 182931 94121 182959
rect 94149 182931 109419 182959
rect 109447 182931 109481 182959
rect 109509 182931 124779 182959
rect 124807 182931 124841 182959
rect 124869 182931 140139 182959
rect 140167 182931 140201 182959
rect 140229 182931 155499 182959
rect 155527 182931 155561 182959
rect 155589 182931 170859 182959
rect 170887 182931 170921 182959
rect 170949 182931 186219 182959
rect 186247 182931 186281 182959
rect 186309 182931 201579 182959
rect 201607 182931 201641 182959
rect 201669 182931 216939 182959
rect 216967 182931 217001 182959
rect 217029 182931 232299 182959
rect 232327 182931 232361 182959
rect 232389 182931 247659 182959
rect 247687 182931 247721 182959
rect 247749 182931 254577 182959
rect 254605 182931 254639 182959
rect 254667 182931 254701 182959
rect 254729 182931 254763 182959
rect 254791 182931 263577 182959
rect 263605 182931 263639 182959
rect 263667 182931 263701 182959
rect 263729 182931 263763 182959
rect 263791 182931 272577 182959
rect 272605 182931 272639 182959
rect 272667 182931 272701 182959
rect 272729 182931 272763 182959
rect 272791 182931 281577 182959
rect 281605 182931 281639 182959
rect 281667 182931 281701 182959
rect 281729 182931 281763 182959
rect 281791 182931 290577 182959
rect 290605 182931 290639 182959
rect 290667 182931 290701 182959
rect 290729 182931 290763 182959
rect 290791 182931 299256 182959
rect 299284 182931 299318 182959
rect 299346 182931 299380 182959
rect 299408 182931 299442 182959
rect 299470 182931 299998 182959
rect -6 182897 299998 182931
rect -6 182869 522 182897
rect 550 182869 584 182897
rect 612 182869 646 182897
rect 674 182869 708 182897
rect 736 182869 2577 182897
rect 2605 182869 2639 182897
rect 2667 182869 2701 182897
rect 2729 182869 2763 182897
rect 2791 182869 11577 182897
rect 11605 182869 11639 182897
rect 11667 182869 11701 182897
rect 11729 182869 11763 182897
rect 11791 182869 17259 182897
rect 17287 182869 17321 182897
rect 17349 182869 20577 182897
rect 20605 182869 20639 182897
rect 20667 182869 20701 182897
rect 20729 182869 20763 182897
rect 20791 182869 29577 182897
rect 29605 182869 29639 182897
rect 29667 182869 29701 182897
rect 29729 182869 29763 182897
rect 29791 182869 32619 182897
rect 32647 182869 32681 182897
rect 32709 182869 47979 182897
rect 48007 182869 48041 182897
rect 48069 182869 63339 182897
rect 63367 182869 63401 182897
rect 63429 182869 78699 182897
rect 78727 182869 78761 182897
rect 78789 182869 94059 182897
rect 94087 182869 94121 182897
rect 94149 182869 109419 182897
rect 109447 182869 109481 182897
rect 109509 182869 124779 182897
rect 124807 182869 124841 182897
rect 124869 182869 140139 182897
rect 140167 182869 140201 182897
rect 140229 182869 155499 182897
rect 155527 182869 155561 182897
rect 155589 182869 170859 182897
rect 170887 182869 170921 182897
rect 170949 182869 186219 182897
rect 186247 182869 186281 182897
rect 186309 182869 201579 182897
rect 201607 182869 201641 182897
rect 201669 182869 216939 182897
rect 216967 182869 217001 182897
rect 217029 182869 232299 182897
rect 232327 182869 232361 182897
rect 232389 182869 247659 182897
rect 247687 182869 247721 182897
rect 247749 182869 254577 182897
rect 254605 182869 254639 182897
rect 254667 182869 254701 182897
rect 254729 182869 254763 182897
rect 254791 182869 263577 182897
rect 263605 182869 263639 182897
rect 263667 182869 263701 182897
rect 263729 182869 263763 182897
rect 263791 182869 272577 182897
rect 272605 182869 272639 182897
rect 272667 182869 272701 182897
rect 272729 182869 272763 182897
rect 272791 182869 281577 182897
rect 281605 182869 281639 182897
rect 281667 182869 281701 182897
rect 281729 182869 281763 182897
rect 281791 182869 290577 182897
rect 290605 182869 290639 182897
rect 290667 182869 290701 182897
rect 290729 182869 290763 182897
rect 290791 182869 299256 182897
rect 299284 182869 299318 182897
rect 299346 182869 299380 182897
rect 299408 182869 299442 182897
rect 299470 182869 299998 182897
rect -6 182835 299998 182869
rect -6 182807 522 182835
rect 550 182807 584 182835
rect 612 182807 646 182835
rect 674 182807 708 182835
rect 736 182807 2577 182835
rect 2605 182807 2639 182835
rect 2667 182807 2701 182835
rect 2729 182807 2763 182835
rect 2791 182807 11577 182835
rect 11605 182807 11639 182835
rect 11667 182807 11701 182835
rect 11729 182807 11763 182835
rect 11791 182807 17259 182835
rect 17287 182807 17321 182835
rect 17349 182807 20577 182835
rect 20605 182807 20639 182835
rect 20667 182807 20701 182835
rect 20729 182807 20763 182835
rect 20791 182807 29577 182835
rect 29605 182807 29639 182835
rect 29667 182807 29701 182835
rect 29729 182807 29763 182835
rect 29791 182807 32619 182835
rect 32647 182807 32681 182835
rect 32709 182807 47979 182835
rect 48007 182807 48041 182835
rect 48069 182807 63339 182835
rect 63367 182807 63401 182835
rect 63429 182807 78699 182835
rect 78727 182807 78761 182835
rect 78789 182807 94059 182835
rect 94087 182807 94121 182835
rect 94149 182807 109419 182835
rect 109447 182807 109481 182835
rect 109509 182807 124779 182835
rect 124807 182807 124841 182835
rect 124869 182807 140139 182835
rect 140167 182807 140201 182835
rect 140229 182807 155499 182835
rect 155527 182807 155561 182835
rect 155589 182807 170859 182835
rect 170887 182807 170921 182835
rect 170949 182807 186219 182835
rect 186247 182807 186281 182835
rect 186309 182807 201579 182835
rect 201607 182807 201641 182835
rect 201669 182807 216939 182835
rect 216967 182807 217001 182835
rect 217029 182807 232299 182835
rect 232327 182807 232361 182835
rect 232389 182807 247659 182835
rect 247687 182807 247721 182835
rect 247749 182807 254577 182835
rect 254605 182807 254639 182835
rect 254667 182807 254701 182835
rect 254729 182807 254763 182835
rect 254791 182807 263577 182835
rect 263605 182807 263639 182835
rect 263667 182807 263701 182835
rect 263729 182807 263763 182835
rect 263791 182807 272577 182835
rect 272605 182807 272639 182835
rect 272667 182807 272701 182835
rect 272729 182807 272763 182835
rect 272791 182807 281577 182835
rect 281605 182807 281639 182835
rect 281667 182807 281701 182835
rect 281729 182807 281763 182835
rect 281791 182807 290577 182835
rect 290605 182807 290639 182835
rect 290667 182807 290701 182835
rect 290729 182807 290763 182835
rect 290791 182807 299256 182835
rect 299284 182807 299318 182835
rect 299346 182807 299380 182835
rect 299408 182807 299442 182835
rect 299470 182807 299998 182835
rect -6 182773 299998 182807
rect -6 182745 522 182773
rect 550 182745 584 182773
rect 612 182745 646 182773
rect 674 182745 708 182773
rect 736 182745 2577 182773
rect 2605 182745 2639 182773
rect 2667 182745 2701 182773
rect 2729 182745 2763 182773
rect 2791 182745 11577 182773
rect 11605 182745 11639 182773
rect 11667 182745 11701 182773
rect 11729 182745 11763 182773
rect 11791 182745 17259 182773
rect 17287 182745 17321 182773
rect 17349 182745 20577 182773
rect 20605 182745 20639 182773
rect 20667 182745 20701 182773
rect 20729 182745 20763 182773
rect 20791 182745 29577 182773
rect 29605 182745 29639 182773
rect 29667 182745 29701 182773
rect 29729 182745 29763 182773
rect 29791 182745 32619 182773
rect 32647 182745 32681 182773
rect 32709 182745 47979 182773
rect 48007 182745 48041 182773
rect 48069 182745 63339 182773
rect 63367 182745 63401 182773
rect 63429 182745 78699 182773
rect 78727 182745 78761 182773
rect 78789 182745 94059 182773
rect 94087 182745 94121 182773
rect 94149 182745 109419 182773
rect 109447 182745 109481 182773
rect 109509 182745 124779 182773
rect 124807 182745 124841 182773
rect 124869 182745 140139 182773
rect 140167 182745 140201 182773
rect 140229 182745 155499 182773
rect 155527 182745 155561 182773
rect 155589 182745 170859 182773
rect 170887 182745 170921 182773
rect 170949 182745 186219 182773
rect 186247 182745 186281 182773
rect 186309 182745 201579 182773
rect 201607 182745 201641 182773
rect 201669 182745 216939 182773
rect 216967 182745 217001 182773
rect 217029 182745 232299 182773
rect 232327 182745 232361 182773
rect 232389 182745 247659 182773
rect 247687 182745 247721 182773
rect 247749 182745 254577 182773
rect 254605 182745 254639 182773
rect 254667 182745 254701 182773
rect 254729 182745 254763 182773
rect 254791 182745 263577 182773
rect 263605 182745 263639 182773
rect 263667 182745 263701 182773
rect 263729 182745 263763 182773
rect 263791 182745 272577 182773
rect 272605 182745 272639 182773
rect 272667 182745 272701 182773
rect 272729 182745 272763 182773
rect 272791 182745 281577 182773
rect 281605 182745 281639 182773
rect 281667 182745 281701 182773
rect 281729 182745 281763 182773
rect 281791 182745 290577 182773
rect 290605 182745 290639 182773
rect 290667 182745 290701 182773
rect 290729 182745 290763 182773
rect 290791 182745 299256 182773
rect 299284 182745 299318 182773
rect 299346 182745 299380 182773
rect 299408 182745 299442 182773
rect 299470 182745 299998 182773
rect -6 182697 299998 182745
rect -6 176959 299998 177007
rect -6 176931 42 176959
rect 70 176931 104 176959
rect 132 176931 166 176959
rect 194 176931 228 176959
rect 256 176931 4437 176959
rect 4465 176931 4499 176959
rect 4527 176931 4561 176959
rect 4589 176931 4623 176959
rect 4651 176931 13437 176959
rect 13465 176931 13499 176959
rect 13527 176931 13561 176959
rect 13589 176931 13623 176959
rect 13651 176931 22437 176959
rect 22465 176931 22499 176959
rect 22527 176931 22561 176959
rect 22589 176931 22623 176959
rect 22651 176931 24939 176959
rect 24967 176931 25001 176959
rect 25029 176931 31437 176959
rect 31465 176931 31499 176959
rect 31527 176931 31561 176959
rect 31589 176931 31623 176959
rect 31651 176931 40299 176959
rect 40327 176931 40361 176959
rect 40389 176931 55659 176959
rect 55687 176931 55721 176959
rect 55749 176931 71019 176959
rect 71047 176931 71081 176959
rect 71109 176931 86379 176959
rect 86407 176931 86441 176959
rect 86469 176931 101739 176959
rect 101767 176931 101801 176959
rect 101829 176931 117099 176959
rect 117127 176931 117161 176959
rect 117189 176931 132459 176959
rect 132487 176931 132521 176959
rect 132549 176931 147819 176959
rect 147847 176931 147881 176959
rect 147909 176931 163179 176959
rect 163207 176931 163241 176959
rect 163269 176931 178539 176959
rect 178567 176931 178601 176959
rect 178629 176931 193899 176959
rect 193927 176931 193961 176959
rect 193989 176931 209259 176959
rect 209287 176931 209321 176959
rect 209349 176931 224619 176959
rect 224647 176931 224681 176959
rect 224709 176931 239979 176959
rect 240007 176931 240041 176959
rect 240069 176931 256437 176959
rect 256465 176931 256499 176959
rect 256527 176931 256561 176959
rect 256589 176931 256623 176959
rect 256651 176931 265437 176959
rect 265465 176931 265499 176959
rect 265527 176931 265561 176959
rect 265589 176931 265623 176959
rect 265651 176931 274437 176959
rect 274465 176931 274499 176959
rect 274527 176931 274561 176959
rect 274589 176931 274623 176959
rect 274651 176931 283437 176959
rect 283465 176931 283499 176959
rect 283527 176931 283561 176959
rect 283589 176931 283623 176959
rect 283651 176931 292437 176959
rect 292465 176931 292499 176959
rect 292527 176931 292561 176959
rect 292589 176931 292623 176959
rect 292651 176931 299736 176959
rect 299764 176931 299798 176959
rect 299826 176931 299860 176959
rect 299888 176931 299922 176959
rect 299950 176931 299998 176959
rect -6 176897 299998 176931
rect -6 176869 42 176897
rect 70 176869 104 176897
rect 132 176869 166 176897
rect 194 176869 228 176897
rect 256 176869 4437 176897
rect 4465 176869 4499 176897
rect 4527 176869 4561 176897
rect 4589 176869 4623 176897
rect 4651 176869 13437 176897
rect 13465 176869 13499 176897
rect 13527 176869 13561 176897
rect 13589 176869 13623 176897
rect 13651 176869 22437 176897
rect 22465 176869 22499 176897
rect 22527 176869 22561 176897
rect 22589 176869 22623 176897
rect 22651 176869 24939 176897
rect 24967 176869 25001 176897
rect 25029 176869 31437 176897
rect 31465 176869 31499 176897
rect 31527 176869 31561 176897
rect 31589 176869 31623 176897
rect 31651 176869 40299 176897
rect 40327 176869 40361 176897
rect 40389 176869 55659 176897
rect 55687 176869 55721 176897
rect 55749 176869 71019 176897
rect 71047 176869 71081 176897
rect 71109 176869 86379 176897
rect 86407 176869 86441 176897
rect 86469 176869 101739 176897
rect 101767 176869 101801 176897
rect 101829 176869 117099 176897
rect 117127 176869 117161 176897
rect 117189 176869 132459 176897
rect 132487 176869 132521 176897
rect 132549 176869 147819 176897
rect 147847 176869 147881 176897
rect 147909 176869 163179 176897
rect 163207 176869 163241 176897
rect 163269 176869 178539 176897
rect 178567 176869 178601 176897
rect 178629 176869 193899 176897
rect 193927 176869 193961 176897
rect 193989 176869 209259 176897
rect 209287 176869 209321 176897
rect 209349 176869 224619 176897
rect 224647 176869 224681 176897
rect 224709 176869 239979 176897
rect 240007 176869 240041 176897
rect 240069 176869 256437 176897
rect 256465 176869 256499 176897
rect 256527 176869 256561 176897
rect 256589 176869 256623 176897
rect 256651 176869 265437 176897
rect 265465 176869 265499 176897
rect 265527 176869 265561 176897
rect 265589 176869 265623 176897
rect 265651 176869 274437 176897
rect 274465 176869 274499 176897
rect 274527 176869 274561 176897
rect 274589 176869 274623 176897
rect 274651 176869 283437 176897
rect 283465 176869 283499 176897
rect 283527 176869 283561 176897
rect 283589 176869 283623 176897
rect 283651 176869 292437 176897
rect 292465 176869 292499 176897
rect 292527 176869 292561 176897
rect 292589 176869 292623 176897
rect 292651 176869 299736 176897
rect 299764 176869 299798 176897
rect 299826 176869 299860 176897
rect 299888 176869 299922 176897
rect 299950 176869 299998 176897
rect -6 176835 299998 176869
rect -6 176807 42 176835
rect 70 176807 104 176835
rect 132 176807 166 176835
rect 194 176807 228 176835
rect 256 176807 4437 176835
rect 4465 176807 4499 176835
rect 4527 176807 4561 176835
rect 4589 176807 4623 176835
rect 4651 176807 13437 176835
rect 13465 176807 13499 176835
rect 13527 176807 13561 176835
rect 13589 176807 13623 176835
rect 13651 176807 22437 176835
rect 22465 176807 22499 176835
rect 22527 176807 22561 176835
rect 22589 176807 22623 176835
rect 22651 176807 24939 176835
rect 24967 176807 25001 176835
rect 25029 176807 31437 176835
rect 31465 176807 31499 176835
rect 31527 176807 31561 176835
rect 31589 176807 31623 176835
rect 31651 176807 40299 176835
rect 40327 176807 40361 176835
rect 40389 176807 55659 176835
rect 55687 176807 55721 176835
rect 55749 176807 71019 176835
rect 71047 176807 71081 176835
rect 71109 176807 86379 176835
rect 86407 176807 86441 176835
rect 86469 176807 101739 176835
rect 101767 176807 101801 176835
rect 101829 176807 117099 176835
rect 117127 176807 117161 176835
rect 117189 176807 132459 176835
rect 132487 176807 132521 176835
rect 132549 176807 147819 176835
rect 147847 176807 147881 176835
rect 147909 176807 163179 176835
rect 163207 176807 163241 176835
rect 163269 176807 178539 176835
rect 178567 176807 178601 176835
rect 178629 176807 193899 176835
rect 193927 176807 193961 176835
rect 193989 176807 209259 176835
rect 209287 176807 209321 176835
rect 209349 176807 224619 176835
rect 224647 176807 224681 176835
rect 224709 176807 239979 176835
rect 240007 176807 240041 176835
rect 240069 176807 256437 176835
rect 256465 176807 256499 176835
rect 256527 176807 256561 176835
rect 256589 176807 256623 176835
rect 256651 176807 265437 176835
rect 265465 176807 265499 176835
rect 265527 176807 265561 176835
rect 265589 176807 265623 176835
rect 265651 176807 274437 176835
rect 274465 176807 274499 176835
rect 274527 176807 274561 176835
rect 274589 176807 274623 176835
rect 274651 176807 283437 176835
rect 283465 176807 283499 176835
rect 283527 176807 283561 176835
rect 283589 176807 283623 176835
rect 283651 176807 292437 176835
rect 292465 176807 292499 176835
rect 292527 176807 292561 176835
rect 292589 176807 292623 176835
rect 292651 176807 299736 176835
rect 299764 176807 299798 176835
rect 299826 176807 299860 176835
rect 299888 176807 299922 176835
rect 299950 176807 299998 176835
rect -6 176773 299998 176807
rect -6 176745 42 176773
rect 70 176745 104 176773
rect 132 176745 166 176773
rect 194 176745 228 176773
rect 256 176745 4437 176773
rect 4465 176745 4499 176773
rect 4527 176745 4561 176773
rect 4589 176745 4623 176773
rect 4651 176745 13437 176773
rect 13465 176745 13499 176773
rect 13527 176745 13561 176773
rect 13589 176745 13623 176773
rect 13651 176745 22437 176773
rect 22465 176745 22499 176773
rect 22527 176745 22561 176773
rect 22589 176745 22623 176773
rect 22651 176745 24939 176773
rect 24967 176745 25001 176773
rect 25029 176745 31437 176773
rect 31465 176745 31499 176773
rect 31527 176745 31561 176773
rect 31589 176745 31623 176773
rect 31651 176745 40299 176773
rect 40327 176745 40361 176773
rect 40389 176745 55659 176773
rect 55687 176745 55721 176773
rect 55749 176745 71019 176773
rect 71047 176745 71081 176773
rect 71109 176745 86379 176773
rect 86407 176745 86441 176773
rect 86469 176745 101739 176773
rect 101767 176745 101801 176773
rect 101829 176745 117099 176773
rect 117127 176745 117161 176773
rect 117189 176745 132459 176773
rect 132487 176745 132521 176773
rect 132549 176745 147819 176773
rect 147847 176745 147881 176773
rect 147909 176745 163179 176773
rect 163207 176745 163241 176773
rect 163269 176745 178539 176773
rect 178567 176745 178601 176773
rect 178629 176745 193899 176773
rect 193927 176745 193961 176773
rect 193989 176745 209259 176773
rect 209287 176745 209321 176773
rect 209349 176745 224619 176773
rect 224647 176745 224681 176773
rect 224709 176745 239979 176773
rect 240007 176745 240041 176773
rect 240069 176745 256437 176773
rect 256465 176745 256499 176773
rect 256527 176745 256561 176773
rect 256589 176745 256623 176773
rect 256651 176745 265437 176773
rect 265465 176745 265499 176773
rect 265527 176745 265561 176773
rect 265589 176745 265623 176773
rect 265651 176745 274437 176773
rect 274465 176745 274499 176773
rect 274527 176745 274561 176773
rect 274589 176745 274623 176773
rect 274651 176745 283437 176773
rect 283465 176745 283499 176773
rect 283527 176745 283561 176773
rect 283589 176745 283623 176773
rect 283651 176745 292437 176773
rect 292465 176745 292499 176773
rect 292527 176745 292561 176773
rect 292589 176745 292623 176773
rect 292651 176745 299736 176773
rect 299764 176745 299798 176773
rect 299826 176745 299860 176773
rect 299888 176745 299922 176773
rect 299950 176745 299998 176773
rect -6 176697 299998 176745
rect -6 173959 299998 174007
rect -6 173931 522 173959
rect 550 173931 584 173959
rect 612 173931 646 173959
rect 674 173931 708 173959
rect 736 173931 2577 173959
rect 2605 173931 2639 173959
rect 2667 173931 2701 173959
rect 2729 173931 2763 173959
rect 2791 173931 11577 173959
rect 11605 173931 11639 173959
rect 11667 173931 11701 173959
rect 11729 173931 11763 173959
rect 11791 173931 17259 173959
rect 17287 173931 17321 173959
rect 17349 173931 20577 173959
rect 20605 173931 20639 173959
rect 20667 173931 20701 173959
rect 20729 173931 20763 173959
rect 20791 173931 29577 173959
rect 29605 173931 29639 173959
rect 29667 173931 29701 173959
rect 29729 173931 29763 173959
rect 29791 173931 32619 173959
rect 32647 173931 32681 173959
rect 32709 173931 47979 173959
rect 48007 173931 48041 173959
rect 48069 173931 63339 173959
rect 63367 173931 63401 173959
rect 63429 173931 78699 173959
rect 78727 173931 78761 173959
rect 78789 173931 94059 173959
rect 94087 173931 94121 173959
rect 94149 173931 109419 173959
rect 109447 173931 109481 173959
rect 109509 173931 124779 173959
rect 124807 173931 124841 173959
rect 124869 173931 140139 173959
rect 140167 173931 140201 173959
rect 140229 173931 155499 173959
rect 155527 173931 155561 173959
rect 155589 173931 170859 173959
rect 170887 173931 170921 173959
rect 170949 173931 186219 173959
rect 186247 173931 186281 173959
rect 186309 173931 201579 173959
rect 201607 173931 201641 173959
rect 201669 173931 216939 173959
rect 216967 173931 217001 173959
rect 217029 173931 232299 173959
rect 232327 173931 232361 173959
rect 232389 173931 247659 173959
rect 247687 173931 247721 173959
rect 247749 173931 254577 173959
rect 254605 173931 254639 173959
rect 254667 173931 254701 173959
rect 254729 173931 254763 173959
rect 254791 173931 263577 173959
rect 263605 173931 263639 173959
rect 263667 173931 263701 173959
rect 263729 173931 263763 173959
rect 263791 173931 272577 173959
rect 272605 173931 272639 173959
rect 272667 173931 272701 173959
rect 272729 173931 272763 173959
rect 272791 173931 281577 173959
rect 281605 173931 281639 173959
rect 281667 173931 281701 173959
rect 281729 173931 281763 173959
rect 281791 173931 290577 173959
rect 290605 173931 290639 173959
rect 290667 173931 290701 173959
rect 290729 173931 290763 173959
rect 290791 173931 299256 173959
rect 299284 173931 299318 173959
rect 299346 173931 299380 173959
rect 299408 173931 299442 173959
rect 299470 173931 299998 173959
rect -6 173897 299998 173931
rect -6 173869 522 173897
rect 550 173869 584 173897
rect 612 173869 646 173897
rect 674 173869 708 173897
rect 736 173869 2577 173897
rect 2605 173869 2639 173897
rect 2667 173869 2701 173897
rect 2729 173869 2763 173897
rect 2791 173869 11577 173897
rect 11605 173869 11639 173897
rect 11667 173869 11701 173897
rect 11729 173869 11763 173897
rect 11791 173869 17259 173897
rect 17287 173869 17321 173897
rect 17349 173869 20577 173897
rect 20605 173869 20639 173897
rect 20667 173869 20701 173897
rect 20729 173869 20763 173897
rect 20791 173869 29577 173897
rect 29605 173869 29639 173897
rect 29667 173869 29701 173897
rect 29729 173869 29763 173897
rect 29791 173869 32619 173897
rect 32647 173869 32681 173897
rect 32709 173869 47979 173897
rect 48007 173869 48041 173897
rect 48069 173869 63339 173897
rect 63367 173869 63401 173897
rect 63429 173869 78699 173897
rect 78727 173869 78761 173897
rect 78789 173869 94059 173897
rect 94087 173869 94121 173897
rect 94149 173869 109419 173897
rect 109447 173869 109481 173897
rect 109509 173869 124779 173897
rect 124807 173869 124841 173897
rect 124869 173869 140139 173897
rect 140167 173869 140201 173897
rect 140229 173869 155499 173897
rect 155527 173869 155561 173897
rect 155589 173869 170859 173897
rect 170887 173869 170921 173897
rect 170949 173869 186219 173897
rect 186247 173869 186281 173897
rect 186309 173869 201579 173897
rect 201607 173869 201641 173897
rect 201669 173869 216939 173897
rect 216967 173869 217001 173897
rect 217029 173869 232299 173897
rect 232327 173869 232361 173897
rect 232389 173869 247659 173897
rect 247687 173869 247721 173897
rect 247749 173869 254577 173897
rect 254605 173869 254639 173897
rect 254667 173869 254701 173897
rect 254729 173869 254763 173897
rect 254791 173869 263577 173897
rect 263605 173869 263639 173897
rect 263667 173869 263701 173897
rect 263729 173869 263763 173897
rect 263791 173869 272577 173897
rect 272605 173869 272639 173897
rect 272667 173869 272701 173897
rect 272729 173869 272763 173897
rect 272791 173869 281577 173897
rect 281605 173869 281639 173897
rect 281667 173869 281701 173897
rect 281729 173869 281763 173897
rect 281791 173869 290577 173897
rect 290605 173869 290639 173897
rect 290667 173869 290701 173897
rect 290729 173869 290763 173897
rect 290791 173869 299256 173897
rect 299284 173869 299318 173897
rect 299346 173869 299380 173897
rect 299408 173869 299442 173897
rect 299470 173869 299998 173897
rect -6 173835 299998 173869
rect -6 173807 522 173835
rect 550 173807 584 173835
rect 612 173807 646 173835
rect 674 173807 708 173835
rect 736 173807 2577 173835
rect 2605 173807 2639 173835
rect 2667 173807 2701 173835
rect 2729 173807 2763 173835
rect 2791 173807 11577 173835
rect 11605 173807 11639 173835
rect 11667 173807 11701 173835
rect 11729 173807 11763 173835
rect 11791 173807 17259 173835
rect 17287 173807 17321 173835
rect 17349 173807 20577 173835
rect 20605 173807 20639 173835
rect 20667 173807 20701 173835
rect 20729 173807 20763 173835
rect 20791 173807 29577 173835
rect 29605 173807 29639 173835
rect 29667 173807 29701 173835
rect 29729 173807 29763 173835
rect 29791 173807 32619 173835
rect 32647 173807 32681 173835
rect 32709 173807 47979 173835
rect 48007 173807 48041 173835
rect 48069 173807 63339 173835
rect 63367 173807 63401 173835
rect 63429 173807 78699 173835
rect 78727 173807 78761 173835
rect 78789 173807 94059 173835
rect 94087 173807 94121 173835
rect 94149 173807 109419 173835
rect 109447 173807 109481 173835
rect 109509 173807 124779 173835
rect 124807 173807 124841 173835
rect 124869 173807 140139 173835
rect 140167 173807 140201 173835
rect 140229 173807 155499 173835
rect 155527 173807 155561 173835
rect 155589 173807 170859 173835
rect 170887 173807 170921 173835
rect 170949 173807 186219 173835
rect 186247 173807 186281 173835
rect 186309 173807 201579 173835
rect 201607 173807 201641 173835
rect 201669 173807 216939 173835
rect 216967 173807 217001 173835
rect 217029 173807 232299 173835
rect 232327 173807 232361 173835
rect 232389 173807 247659 173835
rect 247687 173807 247721 173835
rect 247749 173807 254577 173835
rect 254605 173807 254639 173835
rect 254667 173807 254701 173835
rect 254729 173807 254763 173835
rect 254791 173807 263577 173835
rect 263605 173807 263639 173835
rect 263667 173807 263701 173835
rect 263729 173807 263763 173835
rect 263791 173807 272577 173835
rect 272605 173807 272639 173835
rect 272667 173807 272701 173835
rect 272729 173807 272763 173835
rect 272791 173807 281577 173835
rect 281605 173807 281639 173835
rect 281667 173807 281701 173835
rect 281729 173807 281763 173835
rect 281791 173807 290577 173835
rect 290605 173807 290639 173835
rect 290667 173807 290701 173835
rect 290729 173807 290763 173835
rect 290791 173807 299256 173835
rect 299284 173807 299318 173835
rect 299346 173807 299380 173835
rect 299408 173807 299442 173835
rect 299470 173807 299998 173835
rect -6 173773 299998 173807
rect -6 173745 522 173773
rect 550 173745 584 173773
rect 612 173745 646 173773
rect 674 173745 708 173773
rect 736 173745 2577 173773
rect 2605 173745 2639 173773
rect 2667 173745 2701 173773
rect 2729 173745 2763 173773
rect 2791 173745 11577 173773
rect 11605 173745 11639 173773
rect 11667 173745 11701 173773
rect 11729 173745 11763 173773
rect 11791 173745 17259 173773
rect 17287 173745 17321 173773
rect 17349 173745 20577 173773
rect 20605 173745 20639 173773
rect 20667 173745 20701 173773
rect 20729 173745 20763 173773
rect 20791 173745 29577 173773
rect 29605 173745 29639 173773
rect 29667 173745 29701 173773
rect 29729 173745 29763 173773
rect 29791 173745 32619 173773
rect 32647 173745 32681 173773
rect 32709 173745 47979 173773
rect 48007 173745 48041 173773
rect 48069 173745 63339 173773
rect 63367 173745 63401 173773
rect 63429 173745 78699 173773
rect 78727 173745 78761 173773
rect 78789 173745 94059 173773
rect 94087 173745 94121 173773
rect 94149 173745 109419 173773
rect 109447 173745 109481 173773
rect 109509 173745 124779 173773
rect 124807 173745 124841 173773
rect 124869 173745 140139 173773
rect 140167 173745 140201 173773
rect 140229 173745 155499 173773
rect 155527 173745 155561 173773
rect 155589 173745 170859 173773
rect 170887 173745 170921 173773
rect 170949 173745 186219 173773
rect 186247 173745 186281 173773
rect 186309 173745 201579 173773
rect 201607 173745 201641 173773
rect 201669 173745 216939 173773
rect 216967 173745 217001 173773
rect 217029 173745 232299 173773
rect 232327 173745 232361 173773
rect 232389 173745 247659 173773
rect 247687 173745 247721 173773
rect 247749 173745 254577 173773
rect 254605 173745 254639 173773
rect 254667 173745 254701 173773
rect 254729 173745 254763 173773
rect 254791 173745 263577 173773
rect 263605 173745 263639 173773
rect 263667 173745 263701 173773
rect 263729 173745 263763 173773
rect 263791 173745 272577 173773
rect 272605 173745 272639 173773
rect 272667 173745 272701 173773
rect 272729 173745 272763 173773
rect 272791 173745 281577 173773
rect 281605 173745 281639 173773
rect 281667 173745 281701 173773
rect 281729 173745 281763 173773
rect 281791 173745 290577 173773
rect 290605 173745 290639 173773
rect 290667 173745 290701 173773
rect 290729 173745 290763 173773
rect 290791 173745 299256 173773
rect 299284 173745 299318 173773
rect 299346 173745 299380 173773
rect 299408 173745 299442 173773
rect 299470 173745 299998 173773
rect -6 173697 299998 173745
rect -6 167959 299998 168007
rect -6 167931 42 167959
rect 70 167931 104 167959
rect 132 167931 166 167959
rect 194 167931 228 167959
rect 256 167931 4437 167959
rect 4465 167931 4499 167959
rect 4527 167931 4561 167959
rect 4589 167931 4623 167959
rect 4651 167931 13437 167959
rect 13465 167931 13499 167959
rect 13527 167931 13561 167959
rect 13589 167931 13623 167959
rect 13651 167931 22437 167959
rect 22465 167931 22499 167959
rect 22527 167931 22561 167959
rect 22589 167931 22623 167959
rect 22651 167931 24939 167959
rect 24967 167931 25001 167959
rect 25029 167931 31437 167959
rect 31465 167931 31499 167959
rect 31527 167931 31561 167959
rect 31589 167931 31623 167959
rect 31651 167931 40299 167959
rect 40327 167931 40361 167959
rect 40389 167931 55659 167959
rect 55687 167931 55721 167959
rect 55749 167931 71019 167959
rect 71047 167931 71081 167959
rect 71109 167931 86379 167959
rect 86407 167931 86441 167959
rect 86469 167931 101739 167959
rect 101767 167931 101801 167959
rect 101829 167931 117099 167959
rect 117127 167931 117161 167959
rect 117189 167931 132459 167959
rect 132487 167931 132521 167959
rect 132549 167931 147819 167959
rect 147847 167931 147881 167959
rect 147909 167931 163179 167959
rect 163207 167931 163241 167959
rect 163269 167931 178539 167959
rect 178567 167931 178601 167959
rect 178629 167931 193899 167959
rect 193927 167931 193961 167959
rect 193989 167931 209259 167959
rect 209287 167931 209321 167959
rect 209349 167931 224619 167959
rect 224647 167931 224681 167959
rect 224709 167931 239979 167959
rect 240007 167931 240041 167959
rect 240069 167931 256437 167959
rect 256465 167931 256499 167959
rect 256527 167931 256561 167959
rect 256589 167931 256623 167959
rect 256651 167931 265437 167959
rect 265465 167931 265499 167959
rect 265527 167931 265561 167959
rect 265589 167931 265623 167959
rect 265651 167931 274437 167959
rect 274465 167931 274499 167959
rect 274527 167931 274561 167959
rect 274589 167931 274623 167959
rect 274651 167931 283437 167959
rect 283465 167931 283499 167959
rect 283527 167931 283561 167959
rect 283589 167931 283623 167959
rect 283651 167931 292437 167959
rect 292465 167931 292499 167959
rect 292527 167931 292561 167959
rect 292589 167931 292623 167959
rect 292651 167931 299736 167959
rect 299764 167931 299798 167959
rect 299826 167931 299860 167959
rect 299888 167931 299922 167959
rect 299950 167931 299998 167959
rect -6 167897 299998 167931
rect -6 167869 42 167897
rect 70 167869 104 167897
rect 132 167869 166 167897
rect 194 167869 228 167897
rect 256 167869 4437 167897
rect 4465 167869 4499 167897
rect 4527 167869 4561 167897
rect 4589 167869 4623 167897
rect 4651 167869 13437 167897
rect 13465 167869 13499 167897
rect 13527 167869 13561 167897
rect 13589 167869 13623 167897
rect 13651 167869 22437 167897
rect 22465 167869 22499 167897
rect 22527 167869 22561 167897
rect 22589 167869 22623 167897
rect 22651 167869 24939 167897
rect 24967 167869 25001 167897
rect 25029 167869 31437 167897
rect 31465 167869 31499 167897
rect 31527 167869 31561 167897
rect 31589 167869 31623 167897
rect 31651 167869 40299 167897
rect 40327 167869 40361 167897
rect 40389 167869 55659 167897
rect 55687 167869 55721 167897
rect 55749 167869 71019 167897
rect 71047 167869 71081 167897
rect 71109 167869 86379 167897
rect 86407 167869 86441 167897
rect 86469 167869 101739 167897
rect 101767 167869 101801 167897
rect 101829 167869 117099 167897
rect 117127 167869 117161 167897
rect 117189 167869 132459 167897
rect 132487 167869 132521 167897
rect 132549 167869 147819 167897
rect 147847 167869 147881 167897
rect 147909 167869 163179 167897
rect 163207 167869 163241 167897
rect 163269 167869 178539 167897
rect 178567 167869 178601 167897
rect 178629 167869 193899 167897
rect 193927 167869 193961 167897
rect 193989 167869 209259 167897
rect 209287 167869 209321 167897
rect 209349 167869 224619 167897
rect 224647 167869 224681 167897
rect 224709 167869 239979 167897
rect 240007 167869 240041 167897
rect 240069 167869 256437 167897
rect 256465 167869 256499 167897
rect 256527 167869 256561 167897
rect 256589 167869 256623 167897
rect 256651 167869 265437 167897
rect 265465 167869 265499 167897
rect 265527 167869 265561 167897
rect 265589 167869 265623 167897
rect 265651 167869 274437 167897
rect 274465 167869 274499 167897
rect 274527 167869 274561 167897
rect 274589 167869 274623 167897
rect 274651 167869 283437 167897
rect 283465 167869 283499 167897
rect 283527 167869 283561 167897
rect 283589 167869 283623 167897
rect 283651 167869 292437 167897
rect 292465 167869 292499 167897
rect 292527 167869 292561 167897
rect 292589 167869 292623 167897
rect 292651 167869 299736 167897
rect 299764 167869 299798 167897
rect 299826 167869 299860 167897
rect 299888 167869 299922 167897
rect 299950 167869 299998 167897
rect -6 167835 299998 167869
rect -6 167807 42 167835
rect 70 167807 104 167835
rect 132 167807 166 167835
rect 194 167807 228 167835
rect 256 167807 4437 167835
rect 4465 167807 4499 167835
rect 4527 167807 4561 167835
rect 4589 167807 4623 167835
rect 4651 167807 13437 167835
rect 13465 167807 13499 167835
rect 13527 167807 13561 167835
rect 13589 167807 13623 167835
rect 13651 167807 22437 167835
rect 22465 167807 22499 167835
rect 22527 167807 22561 167835
rect 22589 167807 22623 167835
rect 22651 167807 24939 167835
rect 24967 167807 25001 167835
rect 25029 167807 31437 167835
rect 31465 167807 31499 167835
rect 31527 167807 31561 167835
rect 31589 167807 31623 167835
rect 31651 167807 40299 167835
rect 40327 167807 40361 167835
rect 40389 167807 55659 167835
rect 55687 167807 55721 167835
rect 55749 167807 71019 167835
rect 71047 167807 71081 167835
rect 71109 167807 86379 167835
rect 86407 167807 86441 167835
rect 86469 167807 101739 167835
rect 101767 167807 101801 167835
rect 101829 167807 117099 167835
rect 117127 167807 117161 167835
rect 117189 167807 132459 167835
rect 132487 167807 132521 167835
rect 132549 167807 147819 167835
rect 147847 167807 147881 167835
rect 147909 167807 163179 167835
rect 163207 167807 163241 167835
rect 163269 167807 178539 167835
rect 178567 167807 178601 167835
rect 178629 167807 193899 167835
rect 193927 167807 193961 167835
rect 193989 167807 209259 167835
rect 209287 167807 209321 167835
rect 209349 167807 224619 167835
rect 224647 167807 224681 167835
rect 224709 167807 239979 167835
rect 240007 167807 240041 167835
rect 240069 167807 256437 167835
rect 256465 167807 256499 167835
rect 256527 167807 256561 167835
rect 256589 167807 256623 167835
rect 256651 167807 265437 167835
rect 265465 167807 265499 167835
rect 265527 167807 265561 167835
rect 265589 167807 265623 167835
rect 265651 167807 274437 167835
rect 274465 167807 274499 167835
rect 274527 167807 274561 167835
rect 274589 167807 274623 167835
rect 274651 167807 283437 167835
rect 283465 167807 283499 167835
rect 283527 167807 283561 167835
rect 283589 167807 283623 167835
rect 283651 167807 292437 167835
rect 292465 167807 292499 167835
rect 292527 167807 292561 167835
rect 292589 167807 292623 167835
rect 292651 167807 299736 167835
rect 299764 167807 299798 167835
rect 299826 167807 299860 167835
rect 299888 167807 299922 167835
rect 299950 167807 299998 167835
rect -6 167773 299998 167807
rect -6 167745 42 167773
rect 70 167745 104 167773
rect 132 167745 166 167773
rect 194 167745 228 167773
rect 256 167745 4437 167773
rect 4465 167745 4499 167773
rect 4527 167745 4561 167773
rect 4589 167745 4623 167773
rect 4651 167745 13437 167773
rect 13465 167745 13499 167773
rect 13527 167745 13561 167773
rect 13589 167745 13623 167773
rect 13651 167745 22437 167773
rect 22465 167745 22499 167773
rect 22527 167745 22561 167773
rect 22589 167745 22623 167773
rect 22651 167745 24939 167773
rect 24967 167745 25001 167773
rect 25029 167745 31437 167773
rect 31465 167745 31499 167773
rect 31527 167745 31561 167773
rect 31589 167745 31623 167773
rect 31651 167745 40299 167773
rect 40327 167745 40361 167773
rect 40389 167745 55659 167773
rect 55687 167745 55721 167773
rect 55749 167745 71019 167773
rect 71047 167745 71081 167773
rect 71109 167745 86379 167773
rect 86407 167745 86441 167773
rect 86469 167745 101739 167773
rect 101767 167745 101801 167773
rect 101829 167745 117099 167773
rect 117127 167745 117161 167773
rect 117189 167745 132459 167773
rect 132487 167745 132521 167773
rect 132549 167745 147819 167773
rect 147847 167745 147881 167773
rect 147909 167745 163179 167773
rect 163207 167745 163241 167773
rect 163269 167745 178539 167773
rect 178567 167745 178601 167773
rect 178629 167745 193899 167773
rect 193927 167745 193961 167773
rect 193989 167745 209259 167773
rect 209287 167745 209321 167773
rect 209349 167745 224619 167773
rect 224647 167745 224681 167773
rect 224709 167745 239979 167773
rect 240007 167745 240041 167773
rect 240069 167745 256437 167773
rect 256465 167745 256499 167773
rect 256527 167745 256561 167773
rect 256589 167745 256623 167773
rect 256651 167745 265437 167773
rect 265465 167745 265499 167773
rect 265527 167745 265561 167773
rect 265589 167745 265623 167773
rect 265651 167745 274437 167773
rect 274465 167745 274499 167773
rect 274527 167745 274561 167773
rect 274589 167745 274623 167773
rect 274651 167745 283437 167773
rect 283465 167745 283499 167773
rect 283527 167745 283561 167773
rect 283589 167745 283623 167773
rect 283651 167745 292437 167773
rect 292465 167745 292499 167773
rect 292527 167745 292561 167773
rect 292589 167745 292623 167773
rect 292651 167745 299736 167773
rect 299764 167745 299798 167773
rect 299826 167745 299860 167773
rect 299888 167745 299922 167773
rect 299950 167745 299998 167773
rect -6 167697 299998 167745
rect -6 164959 299998 165007
rect -6 164931 522 164959
rect 550 164931 584 164959
rect 612 164931 646 164959
rect 674 164931 708 164959
rect 736 164931 2577 164959
rect 2605 164931 2639 164959
rect 2667 164931 2701 164959
rect 2729 164931 2763 164959
rect 2791 164931 11577 164959
rect 11605 164931 11639 164959
rect 11667 164931 11701 164959
rect 11729 164931 11763 164959
rect 11791 164931 17259 164959
rect 17287 164931 17321 164959
rect 17349 164931 20577 164959
rect 20605 164931 20639 164959
rect 20667 164931 20701 164959
rect 20729 164931 20763 164959
rect 20791 164931 29577 164959
rect 29605 164931 29639 164959
rect 29667 164931 29701 164959
rect 29729 164931 29763 164959
rect 29791 164931 32619 164959
rect 32647 164931 32681 164959
rect 32709 164931 47979 164959
rect 48007 164931 48041 164959
rect 48069 164931 63339 164959
rect 63367 164931 63401 164959
rect 63429 164931 78699 164959
rect 78727 164931 78761 164959
rect 78789 164931 94059 164959
rect 94087 164931 94121 164959
rect 94149 164931 109419 164959
rect 109447 164931 109481 164959
rect 109509 164931 124779 164959
rect 124807 164931 124841 164959
rect 124869 164931 140139 164959
rect 140167 164931 140201 164959
rect 140229 164931 155499 164959
rect 155527 164931 155561 164959
rect 155589 164931 170859 164959
rect 170887 164931 170921 164959
rect 170949 164931 186219 164959
rect 186247 164931 186281 164959
rect 186309 164931 201579 164959
rect 201607 164931 201641 164959
rect 201669 164931 216939 164959
rect 216967 164931 217001 164959
rect 217029 164931 232299 164959
rect 232327 164931 232361 164959
rect 232389 164931 247659 164959
rect 247687 164931 247721 164959
rect 247749 164931 254577 164959
rect 254605 164931 254639 164959
rect 254667 164931 254701 164959
rect 254729 164931 254763 164959
rect 254791 164931 263577 164959
rect 263605 164931 263639 164959
rect 263667 164931 263701 164959
rect 263729 164931 263763 164959
rect 263791 164931 272577 164959
rect 272605 164931 272639 164959
rect 272667 164931 272701 164959
rect 272729 164931 272763 164959
rect 272791 164931 281577 164959
rect 281605 164931 281639 164959
rect 281667 164931 281701 164959
rect 281729 164931 281763 164959
rect 281791 164931 290577 164959
rect 290605 164931 290639 164959
rect 290667 164931 290701 164959
rect 290729 164931 290763 164959
rect 290791 164931 299256 164959
rect 299284 164931 299318 164959
rect 299346 164931 299380 164959
rect 299408 164931 299442 164959
rect 299470 164931 299998 164959
rect -6 164897 299998 164931
rect -6 164869 522 164897
rect 550 164869 584 164897
rect 612 164869 646 164897
rect 674 164869 708 164897
rect 736 164869 2577 164897
rect 2605 164869 2639 164897
rect 2667 164869 2701 164897
rect 2729 164869 2763 164897
rect 2791 164869 11577 164897
rect 11605 164869 11639 164897
rect 11667 164869 11701 164897
rect 11729 164869 11763 164897
rect 11791 164869 17259 164897
rect 17287 164869 17321 164897
rect 17349 164869 20577 164897
rect 20605 164869 20639 164897
rect 20667 164869 20701 164897
rect 20729 164869 20763 164897
rect 20791 164869 29577 164897
rect 29605 164869 29639 164897
rect 29667 164869 29701 164897
rect 29729 164869 29763 164897
rect 29791 164869 32619 164897
rect 32647 164869 32681 164897
rect 32709 164869 47979 164897
rect 48007 164869 48041 164897
rect 48069 164869 63339 164897
rect 63367 164869 63401 164897
rect 63429 164869 78699 164897
rect 78727 164869 78761 164897
rect 78789 164869 94059 164897
rect 94087 164869 94121 164897
rect 94149 164869 109419 164897
rect 109447 164869 109481 164897
rect 109509 164869 124779 164897
rect 124807 164869 124841 164897
rect 124869 164869 140139 164897
rect 140167 164869 140201 164897
rect 140229 164869 155499 164897
rect 155527 164869 155561 164897
rect 155589 164869 170859 164897
rect 170887 164869 170921 164897
rect 170949 164869 186219 164897
rect 186247 164869 186281 164897
rect 186309 164869 201579 164897
rect 201607 164869 201641 164897
rect 201669 164869 216939 164897
rect 216967 164869 217001 164897
rect 217029 164869 232299 164897
rect 232327 164869 232361 164897
rect 232389 164869 247659 164897
rect 247687 164869 247721 164897
rect 247749 164869 254577 164897
rect 254605 164869 254639 164897
rect 254667 164869 254701 164897
rect 254729 164869 254763 164897
rect 254791 164869 263577 164897
rect 263605 164869 263639 164897
rect 263667 164869 263701 164897
rect 263729 164869 263763 164897
rect 263791 164869 272577 164897
rect 272605 164869 272639 164897
rect 272667 164869 272701 164897
rect 272729 164869 272763 164897
rect 272791 164869 281577 164897
rect 281605 164869 281639 164897
rect 281667 164869 281701 164897
rect 281729 164869 281763 164897
rect 281791 164869 290577 164897
rect 290605 164869 290639 164897
rect 290667 164869 290701 164897
rect 290729 164869 290763 164897
rect 290791 164869 299256 164897
rect 299284 164869 299318 164897
rect 299346 164869 299380 164897
rect 299408 164869 299442 164897
rect 299470 164869 299998 164897
rect -6 164835 299998 164869
rect -6 164807 522 164835
rect 550 164807 584 164835
rect 612 164807 646 164835
rect 674 164807 708 164835
rect 736 164807 2577 164835
rect 2605 164807 2639 164835
rect 2667 164807 2701 164835
rect 2729 164807 2763 164835
rect 2791 164807 11577 164835
rect 11605 164807 11639 164835
rect 11667 164807 11701 164835
rect 11729 164807 11763 164835
rect 11791 164807 17259 164835
rect 17287 164807 17321 164835
rect 17349 164807 20577 164835
rect 20605 164807 20639 164835
rect 20667 164807 20701 164835
rect 20729 164807 20763 164835
rect 20791 164807 29577 164835
rect 29605 164807 29639 164835
rect 29667 164807 29701 164835
rect 29729 164807 29763 164835
rect 29791 164807 32619 164835
rect 32647 164807 32681 164835
rect 32709 164807 47979 164835
rect 48007 164807 48041 164835
rect 48069 164807 63339 164835
rect 63367 164807 63401 164835
rect 63429 164807 78699 164835
rect 78727 164807 78761 164835
rect 78789 164807 94059 164835
rect 94087 164807 94121 164835
rect 94149 164807 109419 164835
rect 109447 164807 109481 164835
rect 109509 164807 124779 164835
rect 124807 164807 124841 164835
rect 124869 164807 140139 164835
rect 140167 164807 140201 164835
rect 140229 164807 155499 164835
rect 155527 164807 155561 164835
rect 155589 164807 170859 164835
rect 170887 164807 170921 164835
rect 170949 164807 186219 164835
rect 186247 164807 186281 164835
rect 186309 164807 201579 164835
rect 201607 164807 201641 164835
rect 201669 164807 216939 164835
rect 216967 164807 217001 164835
rect 217029 164807 232299 164835
rect 232327 164807 232361 164835
rect 232389 164807 247659 164835
rect 247687 164807 247721 164835
rect 247749 164807 254577 164835
rect 254605 164807 254639 164835
rect 254667 164807 254701 164835
rect 254729 164807 254763 164835
rect 254791 164807 263577 164835
rect 263605 164807 263639 164835
rect 263667 164807 263701 164835
rect 263729 164807 263763 164835
rect 263791 164807 272577 164835
rect 272605 164807 272639 164835
rect 272667 164807 272701 164835
rect 272729 164807 272763 164835
rect 272791 164807 281577 164835
rect 281605 164807 281639 164835
rect 281667 164807 281701 164835
rect 281729 164807 281763 164835
rect 281791 164807 290577 164835
rect 290605 164807 290639 164835
rect 290667 164807 290701 164835
rect 290729 164807 290763 164835
rect 290791 164807 299256 164835
rect 299284 164807 299318 164835
rect 299346 164807 299380 164835
rect 299408 164807 299442 164835
rect 299470 164807 299998 164835
rect -6 164773 299998 164807
rect -6 164745 522 164773
rect 550 164745 584 164773
rect 612 164745 646 164773
rect 674 164745 708 164773
rect 736 164745 2577 164773
rect 2605 164745 2639 164773
rect 2667 164745 2701 164773
rect 2729 164745 2763 164773
rect 2791 164745 11577 164773
rect 11605 164745 11639 164773
rect 11667 164745 11701 164773
rect 11729 164745 11763 164773
rect 11791 164745 17259 164773
rect 17287 164745 17321 164773
rect 17349 164745 20577 164773
rect 20605 164745 20639 164773
rect 20667 164745 20701 164773
rect 20729 164745 20763 164773
rect 20791 164745 29577 164773
rect 29605 164745 29639 164773
rect 29667 164745 29701 164773
rect 29729 164745 29763 164773
rect 29791 164745 32619 164773
rect 32647 164745 32681 164773
rect 32709 164745 47979 164773
rect 48007 164745 48041 164773
rect 48069 164745 63339 164773
rect 63367 164745 63401 164773
rect 63429 164745 78699 164773
rect 78727 164745 78761 164773
rect 78789 164745 94059 164773
rect 94087 164745 94121 164773
rect 94149 164745 109419 164773
rect 109447 164745 109481 164773
rect 109509 164745 124779 164773
rect 124807 164745 124841 164773
rect 124869 164745 140139 164773
rect 140167 164745 140201 164773
rect 140229 164745 155499 164773
rect 155527 164745 155561 164773
rect 155589 164745 170859 164773
rect 170887 164745 170921 164773
rect 170949 164745 186219 164773
rect 186247 164745 186281 164773
rect 186309 164745 201579 164773
rect 201607 164745 201641 164773
rect 201669 164745 216939 164773
rect 216967 164745 217001 164773
rect 217029 164745 232299 164773
rect 232327 164745 232361 164773
rect 232389 164745 247659 164773
rect 247687 164745 247721 164773
rect 247749 164745 254577 164773
rect 254605 164745 254639 164773
rect 254667 164745 254701 164773
rect 254729 164745 254763 164773
rect 254791 164745 263577 164773
rect 263605 164745 263639 164773
rect 263667 164745 263701 164773
rect 263729 164745 263763 164773
rect 263791 164745 272577 164773
rect 272605 164745 272639 164773
rect 272667 164745 272701 164773
rect 272729 164745 272763 164773
rect 272791 164745 281577 164773
rect 281605 164745 281639 164773
rect 281667 164745 281701 164773
rect 281729 164745 281763 164773
rect 281791 164745 290577 164773
rect 290605 164745 290639 164773
rect 290667 164745 290701 164773
rect 290729 164745 290763 164773
rect 290791 164745 299256 164773
rect 299284 164745 299318 164773
rect 299346 164745 299380 164773
rect 299408 164745 299442 164773
rect 299470 164745 299998 164773
rect -6 164697 299998 164745
rect -6 158959 299998 159007
rect -6 158931 42 158959
rect 70 158931 104 158959
rect 132 158931 166 158959
rect 194 158931 228 158959
rect 256 158931 4437 158959
rect 4465 158931 4499 158959
rect 4527 158931 4561 158959
rect 4589 158931 4623 158959
rect 4651 158931 13437 158959
rect 13465 158931 13499 158959
rect 13527 158931 13561 158959
rect 13589 158931 13623 158959
rect 13651 158931 22437 158959
rect 22465 158931 22499 158959
rect 22527 158931 22561 158959
rect 22589 158931 22623 158959
rect 22651 158931 24939 158959
rect 24967 158931 25001 158959
rect 25029 158931 31437 158959
rect 31465 158931 31499 158959
rect 31527 158931 31561 158959
rect 31589 158931 31623 158959
rect 31651 158931 40299 158959
rect 40327 158931 40361 158959
rect 40389 158931 55659 158959
rect 55687 158931 55721 158959
rect 55749 158931 71019 158959
rect 71047 158931 71081 158959
rect 71109 158931 86379 158959
rect 86407 158931 86441 158959
rect 86469 158931 101739 158959
rect 101767 158931 101801 158959
rect 101829 158931 117099 158959
rect 117127 158931 117161 158959
rect 117189 158931 132459 158959
rect 132487 158931 132521 158959
rect 132549 158931 147819 158959
rect 147847 158931 147881 158959
rect 147909 158931 163179 158959
rect 163207 158931 163241 158959
rect 163269 158931 178539 158959
rect 178567 158931 178601 158959
rect 178629 158931 193899 158959
rect 193927 158931 193961 158959
rect 193989 158931 209259 158959
rect 209287 158931 209321 158959
rect 209349 158931 224619 158959
rect 224647 158931 224681 158959
rect 224709 158931 239979 158959
rect 240007 158931 240041 158959
rect 240069 158931 256437 158959
rect 256465 158931 256499 158959
rect 256527 158931 256561 158959
rect 256589 158931 256623 158959
rect 256651 158931 265437 158959
rect 265465 158931 265499 158959
rect 265527 158931 265561 158959
rect 265589 158931 265623 158959
rect 265651 158931 274437 158959
rect 274465 158931 274499 158959
rect 274527 158931 274561 158959
rect 274589 158931 274623 158959
rect 274651 158931 283437 158959
rect 283465 158931 283499 158959
rect 283527 158931 283561 158959
rect 283589 158931 283623 158959
rect 283651 158931 292437 158959
rect 292465 158931 292499 158959
rect 292527 158931 292561 158959
rect 292589 158931 292623 158959
rect 292651 158931 299736 158959
rect 299764 158931 299798 158959
rect 299826 158931 299860 158959
rect 299888 158931 299922 158959
rect 299950 158931 299998 158959
rect -6 158897 299998 158931
rect -6 158869 42 158897
rect 70 158869 104 158897
rect 132 158869 166 158897
rect 194 158869 228 158897
rect 256 158869 4437 158897
rect 4465 158869 4499 158897
rect 4527 158869 4561 158897
rect 4589 158869 4623 158897
rect 4651 158869 13437 158897
rect 13465 158869 13499 158897
rect 13527 158869 13561 158897
rect 13589 158869 13623 158897
rect 13651 158869 22437 158897
rect 22465 158869 22499 158897
rect 22527 158869 22561 158897
rect 22589 158869 22623 158897
rect 22651 158869 24939 158897
rect 24967 158869 25001 158897
rect 25029 158869 31437 158897
rect 31465 158869 31499 158897
rect 31527 158869 31561 158897
rect 31589 158869 31623 158897
rect 31651 158869 40299 158897
rect 40327 158869 40361 158897
rect 40389 158869 55659 158897
rect 55687 158869 55721 158897
rect 55749 158869 71019 158897
rect 71047 158869 71081 158897
rect 71109 158869 86379 158897
rect 86407 158869 86441 158897
rect 86469 158869 101739 158897
rect 101767 158869 101801 158897
rect 101829 158869 117099 158897
rect 117127 158869 117161 158897
rect 117189 158869 132459 158897
rect 132487 158869 132521 158897
rect 132549 158869 147819 158897
rect 147847 158869 147881 158897
rect 147909 158869 163179 158897
rect 163207 158869 163241 158897
rect 163269 158869 178539 158897
rect 178567 158869 178601 158897
rect 178629 158869 193899 158897
rect 193927 158869 193961 158897
rect 193989 158869 209259 158897
rect 209287 158869 209321 158897
rect 209349 158869 224619 158897
rect 224647 158869 224681 158897
rect 224709 158869 239979 158897
rect 240007 158869 240041 158897
rect 240069 158869 256437 158897
rect 256465 158869 256499 158897
rect 256527 158869 256561 158897
rect 256589 158869 256623 158897
rect 256651 158869 265437 158897
rect 265465 158869 265499 158897
rect 265527 158869 265561 158897
rect 265589 158869 265623 158897
rect 265651 158869 274437 158897
rect 274465 158869 274499 158897
rect 274527 158869 274561 158897
rect 274589 158869 274623 158897
rect 274651 158869 283437 158897
rect 283465 158869 283499 158897
rect 283527 158869 283561 158897
rect 283589 158869 283623 158897
rect 283651 158869 292437 158897
rect 292465 158869 292499 158897
rect 292527 158869 292561 158897
rect 292589 158869 292623 158897
rect 292651 158869 299736 158897
rect 299764 158869 299798 158897
rect 299826 158869 299860 158897
rect 299888 158869 299922 158897
rect 299950 158869 299998 158897
rect -6 158835 299998 158869
rect -6 158807 42 158835
rect 70 158807 104 158835
rect 132 158807 166 158835
rect 194 158807 228 158835
rect 256 158807 4437 158835
rect 4465 158807 4499 158835
rect 4527 158807 4561 158835
rect 4589 158807 4623 158835
rect 4651 158807 13437 158835
rect 13465 158807 13499 158835
rect 13527 158807 13561 158835
rect 13589 158807 13623 158835
rect 13651 158807 22437 158835
rect 22465 158807 22499 158835
rect 22527 158807 22561 158835
rect 22589 158807 22623 158835
rect 22651 158807 24939 158835
rect 24967 158807 25001 158835
rect 25029 158807 31437 158835
rect 31465 158807 31499 158835
rect 31527 158807 31561 158835
rect 31589 158807 31623 158835
rect 31651 158807 40299 158835
rect 40327 158807 40361 158835
rect 40389 158807 55659 158835
rect 55687 158807 55721 158835
rect 55749 158807 71019 158835
rect 71047 158807 71081 158835
rect 71109 158807 86379 158835
rect 86407 158807 86441 158835
rect 86469 158807 101739 158835
rect 101767 158807 101801 158835
rect 101829 158807 117099 158835
rect 117127 158807 117161 158835
rect 117189 158807 132459 158835
rect 132487 158807 132521 158835
rect 132549 158807 147819 158835
rect 147847 158807 147881 158835
rect 147909 158807 163179 158835
rect 163207 158807 163241 158835
rect 163269 158807 178539 158835
rect 178567 158807 178601 158835
rect 178629 158807 193899 158835
rect 193927 158807 193961 158835
rect 193989 158807 209259 158835
rect 209287 158807 209321 158835
rect 209349 158807 224619 158835
rect 224647 158807 224681 158835
rect 224709 158807 239979 158835
rect 240007 158807 240041 158835
rect 240069 158807 256437 158835
rect 256465 158807 256499 158835
rect 256527 158807 256561 158835
rect 256589 158807 256623 158835
rect 256651 158807 265437 158835
rect 265465 158807 265499 158835
rect 265527 158807 265561 158835
rect 265589 158807 265623 158835
rect 265651 158807 274437 158835
rect 274465 158807 274499 158835
rect 274527 158807 274561 158835
rect 274589 158807 274623 158835
rect 274651 158807 283437 158835
rect 283465 158807 283499 158835
rect 283527 158807 283561 158835
rect 283589 158807 283623 158835
rect 283651 158807 292437 158835
rect 292465 158807 292499 158835
rect 292527 158807 292561 158835
rect 292589 158807 292623 158835
rect 292651 158807 299736 158835
rect 299764 158807 299798 158835
rect 299826 158807 299860 158835
rect 299888 158807 299922 158835
rect 299950 158807 299998 158835
rect -6 158773 299998 158807
rect -6 158745 42 158773
rect 70 158745 104 158773
rect 132 158745 166 158773
rect 194 158745 228 158773
rect 256 158745 4437 158773
rect 4465 158745 4499 158773
rect 4527 158745 4561 158773
rect 4589 158745 4623 158773
rect 4651 158745 13437 158773
rect 13465 158745 13499 158773
rect 13527 158745 13561 158773
rect 13589 158745 13623 158773
rect 13651 158745 22437 158773
rect 22465 158745 22499 158773
rect 22527 158745 22561 158773
rect 22589 158745 22623 158773
rect 22651 158745 24939 158773
rect 24967 158745 25001 158773
rect 25029 158745 31437 158773
rect 31465 158745 31499 158773
rect 31527 158745 31561 158773
rect 31589 158745 31623 158773
rect 31651 158745 40299 158773
rect 40327 158745 40361 158773
rect 40389 158745 55659 158773
rect 55687 158745 55721 158773
rect 55749 158745 71019 158773
rect 71047 158745 71081 158773
rect 71109 158745 86379 158773
rect 86407 158745 86441 158773
rect 86469 158745 101739 158773
rect 101767 158745 101801 158773
rect 101829 158745 117099 158773
rect 117127 158745 117161 158773
rect 117189 158745 132459 158773
rect 132487 158745 132521 158773
rect 132549 158745 147819 158773
rect 147847 158745 147881 158773
rect 147909 158745 163179 158773
rect 163207 158745 163241 158773
rect 163269 158745 178539 158773
rect 178567 158745 178601 158773
rect 178629 158745 193899 158773
rect 193927 158745 193961 158773
rect 193989 158745 209259 158773
rect 209287 158745 209321 158773
rect 209349 158745 224619 158773
rect 224647 158745 224681 158773
rect 224709 158745 239979 158773
rect 240007 158745 240041 158773
rect 240069 158745 256437 158773
rect 256465 158745 256499 158773
rect 256527 158745 256561 158773
rect 256589 158745 256623 158773
rect 256651 158745 265437 158773
rect 265465 158745 265499 158773
rect 265527 158745 265561 158773
rect 265589 158745 265623 158773
rect 265651 158745 274437 158773
rect 274465 158745 274499 158773
rect 274527 158745 274561 158773
rect 274589 158745 274623 158773
rect 274651 158745 283437 158773
rect 283465 158745 283499 158773
rect 283527 158745 283561 158773
rect 283589 158745 283623 158773
rect 283651 158745 292437 158773
rect 292465 158745 292499 158773
rect 292527 158745 292561 158773
rect 292589 158745 292623 158773
rect 292651 158745 299736 158773
rect 299764 158745 299798 158773
rect 299826 158745 299860 158773
rect 299888 158745 299922 158773
rect 299950 158745 299998 158773
rect -6 158697 299998 158745
rect -6 155959 299998 156007
rect -6 155931 522 155959
rect 550 155931 584 155959
rect 612 155931 646 155959
rect 674 155931 708 155959
rect 736 155931 2577 155959
rect 2605 155931 2639 155959
rect 2667 155931 2701 155959
rect 2729 155931 2763 155959
rect 2791 155931 11577 155959
rect 11605 155931 11639 155959
rect 11667 155931 11701 155959
rect 11729 155931 11763 155959
rect 11791 155931 17259 155959
rect 17287 155931 17321 155959
rect 17349 155931 20577 155959
rect 20605 155931 20639 155959
rect 20667 155931 20701 155959
rect 20729 155931 20763 155959
rect 20791 155931 29577 155959
rect 29605 155931 29639 155959
rect 29667 155931 29701 155959
rect 29729 155931 29763 155959
rect 29791 155931 32619 155959
rect 32647 155931 32681 155959
rect 32709 155931 47979 155959
rect 48007 155931 48041 155959
rect 48069 155931 63339 155959
rect 63367 155931 63401 155959
rect 63429 155931 78699 155959
rect 78727 155931 78761 155959
rect 78789 155931 94059 155959
rect 94087 155931 94121 155959
rect 94149 155931 109419 155959
rect 109447 155931 109481 155959
rect 109509 155931 124779 155959
rect 124807 155931 124841 155959
rect 124869 155931 140139 155959
rect 140167 155931 140201 155959
rect 140229 155931 155499 155959
rect 155527 155931 155561 155959
rect 155589 155931 170859 155959
rect 170887 155931 170921 155959
rect 170949 155931 186219 155959
rect 186247 155931 186281 155959
rect 186309 155931 201579 155959
rect 201607 155931 201641 155959
rect 201669 155931 216939 155959
rect 216967 155931 217001 155959
rect 217029 155931 232299 155959
rect 232327 155931 232361 155959
rect 232389 155931 247659 155959
rect 247687 155931 247721 155959
rect 247749 155931 254577 155959
rect 254605 155931 254639 155959
rect 254667 155931 254701 155959
rect 254729 155931 254763 155959
rect 254791 155931 263577 155959
rect 263605 155931 263639 155959
rect 263667 155931 263701 155959
rect 263729 155931 263763 155959
rect 263791 155931 272577 155959
rect 272605 155931 272639 155959
rect 272667 155931 272701 155959
rect 272729 155931 272763 155959
rect 272791 155931 281577 155959
rect 281605 155931 281639 155959
rect 281667 155931 281701 155959
rect 281729 155931 281763 155959
rect 281791 155931 290577 155959
rect 290605 155931 290639 155959
rect 290667 155931 290701 155959
rect 290729 155931 290763 155959
rect 290791 155931 299256 155959
rect 299284 155931 299318 155959
rect 299346 155931 299380 155959
rect 299408 155931 299442 155959
rect 299470 155931 299998 155959
rect -6 155897 299998 155931
rect -6 155869 522 155897
rect 550 155869 584 155897
rect 612 155869 646 155897
rect 674 155869 708 155897
rect 736 155869 2577 155897
rect 2605 155869 2639 155897
rect 2667 155869 2701 155897
rect 2729 155869 2763 155897
rect 2791 155869 11577 155897
rect 11605 155869 11639 155897
rect 11667 155869 11701 155897
rect 11729 155869 11763 155897
rect 11791 155869 17259 155897
rect 17287 155869 17321 155897
rect 17349 155869 20577 155897
rect 20605 155869 20639 155897
rect 20667 155869 20701 155897
rect 20729 155869 20763 155897
rect 20791 155869 29577 155897
rect 29605 155869 29639 155897
rect 29667 155869 29701 155897
rect 29729 155869 29763 155897
rect 29791 155869 32619 155897
rect 32647 155869 32681 155897
rect 32709 155869 47979 155897
rect 48007 155869 48041 155897
rect 48069 155869 63339 155897
rect 63367 155869 63401 155897
rect 63429 155869 78699 155897
rect 78727 155869 78761 155897
rect 78789 155869 94059 155897
rect 94087 155869 94121 155897
rect 94149 155869 109419 155897
rect 109447 155869 109481 155897
rect 109509 155869 124779 155897
rect 124807 155869 124841 155897
rect 124869 155869 140139 155897
rect 140167 155869 140201 155897
rect 140229 155869 155499 155897
rect 155527 155869 155561 155897
rect 155589 155869 170859 155897
rect 170887 155869 170921 155897
rect 170949 155869 186219 155897
rect 186247 155869 186281 155897
rect 186309 155869 201579 155897
rect 201607 155869 201641 155897
rect 201669 155869 216939 155897
rect 216967 155869 217001 155897
rect 217029 155869 232299 155897
rect 232327 155869 232361 155897
rect 232389 155869 247659 155897
rect 247687 155869 247721 155897
rect 247749 155869 254577 155897
rect 254605 155869 254639 155897
rect 254667 155869 254701 155897
rect 254729 155869 254763 155897
rect 254791 155869 263577 155897
rect 263605 155869 263639 155897
rect 263667 155869 263701 155897
rect 263729 155869 263763 155897
rect 263791 155869 272577 155897
rect 272605 155869 272639 155897
rect 272667 155869 272701 155897
rect 272729 155869 272763 155897
rect 272791 155869 281577 155897
rect 281605 155869 281639 155897
rect 281667 155869 281701 155897
rect 281729 155869 281763 155897
rect 281791 155869 290577 155897
rect 290605 155869 290639 155897
rect 290667 155869 290701 155897
rect 290729 155869 290763 155897
rect 290791 155869 299256 155897
rect 299284 155869 299318 155897
rect 299346 155869 299380 155897
rect 299408 155869 299442 155897
rect 299470 155869 299998 155897
rect -6 155835 299998 155869
rect -6 155807 522 155835
rect 550 155807 584 155835
rect 612 155807 646 155835
rect 674 155807 708 155835
rect 736 155807 2577 155835
rect 2605 155807 2639 155835
rect 2667 155807 2701 155835
rect 2729 155807 2763 155835
rect 2791 155807 11577 155835
rect 11605 155807 11639 155835
rect 11667 155807 11701 155835
rect 11729 155807 11763 155835
rect 11791 155807 17259 155835
rect 17287 155807 17321 155835
rect 17349 155807 20577 155835
rect 20605 155807 20639 155835
rect 20667 155807 20701 155835
rect 20729 155807 20763 155835
rect 20791 155807 29577 155835
rect 29605 155807 29639 155835
rect 29667 155807 29701 155835
rect 29729 155807 29763 155835
rect 29791 155807 32619 155835
rect 32647 155807 32681 155835
rect 32709 155807 47979 155835
rect 48007 155807 48041 155835
rect 48069 155807 63339 155835
rect 63367 155807 63401 155835
rect 63429 155807 78699 155835
rect 78727 155807 78761 155835
rect 78789 155807 94059 155835
rect 94087 155807 94121 155835
rect 94149 155807 109419 155835
rect 109447 155807 109481 155835
rect 109509 155807 124779 155835
rect 124807 155807 124841 155835
rect 124869 155807 140139 155835
rect 140167 155807 140201 155835
rect 140229 155807 155499 155835
rect 155527 155807 155561 155835
rect 155589 155807 170859 155835
rect 170887 155807 170921 155835
rect 170949 155807 186219 155835
rect 186247 155807 186281 155835
rect 186309 155807 201579 155835
rect 201607 155807 201641 155835
rect 201669 155807 216939 155835
rect 216967 155807 217001 155835
rect 217029 155807 232299 155835
rect 232327 155807 232361 155835
rect 232389 155807 247659 155835
rect 247687 155807 247721 155835
rect 247749 155807 254577 155835
rect 254605 155807 254639 155835
rect 254667 155807 254701 155835
rect 254729 155807 254763 155835
rect 254791 155807 263577 155835
rect 263605 155807 263639 155835
rect 263667 155807 263701 155835
rect 263729 155807 263763 155835
rect 263791 155807 272577 155835
rect 272605 155807 272639 155835
rect 272667 155807 272701 155835
rect 272729 155807 272763 155835
rect 272791 155807 281577 155835
rect 281605 155807 281639 155835
rect 281667 155807 281701 155835
rect 281729 155807 281763 155835
rect 281791 155807 290577 155835
rect 290605 155807 290639 155835
rect 290667 155807 290701 155835
rect 290729 155807 290763 155835
rect 290791 155807 299256 155835
rect 299284 155807 299318 155835
rect 299346 155807 299380 155835
rect 299408 155807 299442 155835
rect 299470 155807 299998 155835
rect -6 155773 299998 155807
rect -6 155745 522 155773
rect 550 155745 584 155773
rect 612 155745 646 155773
rect 674 155745 708 155773
rect 736 155745 2577 155773
rect 2605 155745 2639 155773
rect 2667 155745 2701 155773
rect 2729 155745 2763 155773
rect 2791 155745 11577 155773
rect 11605 155745 11639 155773
rect 11667 155745 11701 155773
rect 11729 155745 11763 155773
rect 11791 155745 17259 155773
rect 17287 155745 17321 155773
rect 17349 155745 20577 155773
rect 20605 155745 20639 155773
rect 20667 155745 20701 155773
rect 20729 155745 20763 155773
rect 20791 155745 29577 155773
rect 29605 155745 29639 155773
rect 29667 155745 29701 155773
rect 29729 155745 29763 155773
rect 29791 155745 32619 155773
rect 32647 155745 32681 155773
rect 32709 155745 47979 155773
rect 48007 155745 48041 155773
rect 48069 155745 63339 155773
rect 63367 155745 63401 155773
rect 63429 155745 78699 155773
rect 78727 155745 78761 155773
rect 78789 155745 94059 155773
rect 94087 155745 94121 155773
rect 94149 155745 109419 155773
rect 109447 155745 109481 155773
rect 109509 155745 124779 155773
rect 124807 155745 124841 155773
rect 124869 155745 140139 155773
rect 140167 155745 140201 155773
rect 140229 155745 155499 155773
rect 155527 155745 155561 155773
rect 155589 155745 170859 155773
rect 170887 155745 170921 155773
rect 170949 155745 186219 155773
rect 186247 155745 186281 155773
rect 186309 155745 201579 155773
rect 201607 155745 201641 155773
rect 201669 155745 216939 155773
rect 216967 155745 217001 155773
rect 217029 155745 232299 155773
rect 232327 155745 232361 155773
rect 232389 155745 247659 155773
rect 247687 155745 247721 155773
rect 247749 155745 254577 155773
rect 254605 155745 254639 155773
rect 254667 155745 254701 155773
rect 254729 155745 254763 155773
rect 254791 155745 263577 155773
rect 263605 155745 263639 155773
rect 263667 155745 263701 155773
rect 263729 155745 263763 155773
rect 263791 155745 272577 155773
rect 272605 155745 272639 155773
rect 272667 155745 272701 155773
rect 272729 155745 272763 155773
rect 272791 155745 281577 155773
rect 281605 155745 281639 155773
rect 281667 155745 281701 155773
rect 281729 155745 281763 155773
rect 281791 155745 290577 155773
rect 290605 155745 290639 155773
rect 290667 155745 290701 155773
rect 290729 155745 290763 155773
rect 290791 155745 299256 155773
rect 299284 155745 299318 155773
rect 299346 155745 299380 155773
rect 299408 155745 299442 155773
rect 299470 155745 299998 155773
rect -6 155697 299998 155745
rect -6 149959 299998 150007
rect -6 149931 42 149959
rect 70 149931 104 149959
rect 132 149931 166 149959
rect 194 149931 228 149959
rect 256 149931 4437 149959
rect 4465 149931 4499 149959
rect 4527 149931 4561 149959
rect 4589 149931 4623 149959
rect 4651 149931 13437 149959
rect 13465 149931 13499 149959
rect 13527 149931 13561 149959
rect 13589 149931 13623 149959
rect 13651 149931 22437 149959
rect 22465 149931 22499 149959
rect 22527 149931 22561 149959
rect 22589 149931 22623 149959
rect 22651 149931 24939 149959
rect 24967 149931 25001 149959
rect 25029 149931 31437 149959
rect 31465 149931 31499 149959
rect 31527 149931 31561 149959
rect 31589 149931 31623 149959
rect 31651 149931 40299 149959
rect 40327 149931 40361 149959
rect 40389 149931 55659 149959
rect 55687 149931 55721 149959
rect 55749 149931 71019 149959
rect 71047 149931 71081 149959
rect 71109 149931 86379 149959
rect 86407 149931 86441 149959
rect 86469 149931 101739 149959
rect 101767 149931 101801 149959
rect 101829 149931 117099 149959
rect 117127 149931 117161 149959
rect 117189 149931 132459 149959
rect 132487 149931 132521 149959
rect 132549 149931 147819 149959
rect 147847 149931 147881 149959
rect 147909 149931 163179 149959
rect 163207 149931 163241 149959
rect 163269 149931 178539 149959
rect 178567 149931 178601 149959
rect 178629 149931 193899 149959
rect 193927 149931 193961 149959
rect 193989 149931 209259 149959
rect 209287 149931 209321 149959
rect 209349 149931 224619 149959
rect 224647 149931 224681 149959
rect 224709 149931 239979 149959
rect 240007 149931 240041 149959
rect 240069 149931 256437 149959
rect 256465 149931 256499 149959
rect 256527 149931 256561 149959
rect 256589 149931 256623 149959
rect 256651 149931 265437 149959
rect 265465 149931 265499 149959
rect 265527 149931 265561 149959
rect 265589 149931 265623 149959
rect 265651 149931 274437 149959
rect 274465 149931 274499 149959
rect 274527 149931 274561 149959
rect 274589 149931 274623 149959
rect 274651 149931 283437 149959
rect 283465 149931 283499 149959
rect 283527 149931 283561 149959
rect 283589 149931 283623 149959
rect 283651 149931 292437 149959
rect 292465 149931 292499 149959
rect 292527 149931 292561 149959
rect 292589 149931 292623 149959
rect 292651 149931 299736 149959
rect 299764 149931 299798 149959
rect 299826 149931 299860 149959
rect 299888 149931 299922 149959
rect 299950 149931 299998 149959
rect -6 149897 299998 149931
rect -6 149869 42 149897
rect 70 149869 104 149897
rect 132 149869 166 149897
rect 194 149869 228 149897
rect 256 149869 4437 149897
rect 4465 149869 4499 149897
rect 4527 149869 4561 149897
rect 4589 149869 4623 149897
rect 4651 149869 13437 149897
rect 13465 149869 13499 149897
rect 13527 149869 13561 149897
rect 13589 149869 13623 149897
rect 13651 149869 22437 149897
rect 22465 149869 22499 149897
rect 22527 149869 22561 149897
rect 22589 149869 22623 149897
rect 22651 149869 24939 149897
rect 24967 149869 25001 149897
rect 25029 149869 31437 149897
rect 31465 149869 31499 149897
rect 31527 149869 31561 149897
rect 31589 149869 31623 149897
rect 31651 149869 40299 149897
rect 40327 149869 40361 149897
rect 40389 149869 55659 149897
rect 55687 149869 55721 149897
rect 55749 149869 71019 149897
rect 71047 149869 71081 149897
rect 71109 149869 86379 149897
rect 86407 149869 86441 149897
rect 86469 149869 101739 149897
rect 101767 149869 101801 149897
rect 101829 149869 117099 149897
rect 117127 149869 117161 149897
rect 117189 149869 132459 149897
rect 132487 149869 132521 149897
rect 132549 149869 147819 149897
rect 147847 149869 147881 149897
rect 147909 149869 163179 149897
rect 163207 149869 163241 149897
rect 163269 149869 178539 149897
rect 178567 149869 178601 149897
rect 178629 149869 193899 149897
rect 193927 149869 193961 149897
rect 193989 149869 209259 149897
rect 209287 149869 209321 149897
rect 209349 149869 224619 149897
rect 224647 149869 224681 149897
rect 224709 149869 239979 149897
rect 240007 149869 240041 149897
rect 240069 149869 256437 149897
rect 256465 149869 256499 149897
rect 256527 149869 256561 149897
rect 256589 149869 256623 149897
rect 256651 149869 265437 149897
rect 265465 149869 265499 149897
rect 265527 149869 265561 149897
rect 265589 149869 265623 149897
rect 265651 149869 274437 149897
rect 274465 149869 274499 149897
rect 274527 149869 274561 149897
rect 274589 149869 274623 149897
rect 274651 149869 283437 149897
rect 283465 149869 283499 149897
rect 283527 149869 283561 149897
rect 283589 149869 283623 149897
rect 283651 149869 292437 149897
rect 292465 149869 292499 149897
rect 292527 149869 292561 149897
rect 292589 149869 292623 149897
rect 292651 149869 299736 149897
rect 299764 149869 299798 149897
rect 299826 149869 299860 149897
rect 299888 149869 299922 149897
rect 299950 149869 299998 149897
rect -6 149835 299998 149869
rect -6 149807 42 149835
rect 70 149807 104 149835
rect 132 149807 166 149835
rect 194 149807 228 149835
rect 256 149807 4437 149835
rect 4465 149807 4499 149835
rect 4527 149807 4561 149835
rect 4589 149807 4623 149835
rect 4651 149807 13437 149835
rect 13465 149807 13499 149835
rect 13527 149807 13561 149835
rect 13589 149807 13623 149835
rect 13651 149807 22437 149835
rect 22465 149807 22499 149835
rect 22527 149807 22561 149835
rect 22589 149807 22623 149835
rect 22651 149807 24939 149835
rect 24967 149807 25001 149835
rect 25029 149807 31437 149835
rect 31465 149807 31499 149835
rect 31527 149807 31561 149835
rect 31589 149807 31623 149835
rect 31651 149807 40299 149835
rect 40327 149807 40361 149835
rect 40389 149807 55659 149835
rect 55687 149807 55721 149835
rect 55749 149807 71019 149835
rect 71047 149807 71081 149835
rect 71109 149807 86379 149835
rect 86407 149807 86441 149835
rect 86469 149807 101739 149835
rect 101767 149807 101801 149835
rect 101829 149807 117099 149835
rect 117127 149807 117161 149835
rect 117189 149807 132459 149835
rect 132487 149807 132521 149835
rect 132549 149807 147819 149835
rect 147847 149807 147881 149835
rect 147909 149807 163179 149835
rect 163207 149807 163241 149835
rect 163269 149807 178539 149835
rect 178567 149807 178601 149835
rect 178629 149807 193899 149835
rect 193927 149807 193961 149835
rect 193989 149807 209259 149835
rect 209287 149807 209321 149835
rect 209349 149807 224619 149835
rect 224647 149807 224681 149835
rect 224709 149807 239979 149835
rect 240007 149807 240041 149835
rect 240069 149807 256437 149835
rect 256465 149807 256499 149835
rect 256527 149807 256561 149835
rect 256589 149807 256623 149835
rect 256651 149807 265437 149835
rect 265465 149807 265499 149835
rect 265527 149807 265561 149835
rect 265589 149807 265623 149835
rect 265651 149807 274437 149835
rect 274465 149807 274499 149835
rect 274527 149807 274561 149835
rect 274589 149807 274623 149835
rect 274651 149807 283437 149835
rect 283465 149807 283499 149835
rect 283527 149807 283561 149835
rect 283589 149807 283623 149835
rect 283651 149807 292437 149835
rect 292465 149807 292499 149835
rect 292527 149807 292561 149835
rect 292589 149807 292623 149835
rect 292651 149807 299736 149835
rect 299764 149807 299798 149835
rect 299826 149807 299860 149835
rect 299888 149807 299922 149835
rect 299950 149807 299998 149835
rect -6 149773 299998 149807
rect -6 149745 42 149773
rect 70 149745 104 149773
rect 132 149745 166 149773
rect 194 149745 228 149773
rect 256 149745 4437 149773
rect 4465 149745 4499 149773
rect 4527 149745 4561 149773
rect 4589 149745 4623 149773
rect 4651 149745 13437 149773
rect 13465 149745 13499 149773
rect 13527 149745 13561 149773
rect 13589 149745 13623 149773
rect 13651 149745 22437 149773
rect 22465 149745 22499 149773
rect 22527 149745 22561 149773
rect 22589 149745 22623 149773
rect 22651 149745 24939 149773
rect 24967 149745 25001 149773
rect 25029 149745 31437 149773
rect 31465 149745 31499 149773
rect 31527 149745 31561 149773
rect 31589 149745 31623 149773
rect 31651 149745 40299 149773
rect 40327 149745 40361 149773
rect 40389 149745 55659 149773
rect 55687 149745 55721 149773
rect 55749 149745 71019 149773
rect 71047 149745 71081 149773
rect 71109 149745 86379 149773
rect 86407 149745 86441 149773
rect 86469 149745 101739 149773
rect 101767 149745 101801 149773
rect 101829 149745 117099 149773
rect 117127 149745 117161 149773
rect 117189 149745 132459 149773
rect 132487 149745 132521 149773
rect 132549 149745 147819 149773
rect 147847 149745 147881 149773
rect 147909 149745 163179 149773
rect 163207 149745 163241 149773
rect 163269 149745 178539 149773
rect 178567 149745 178601 149773
rect 178629 149745 193899 149773
rect 193927 149745 193961 149773
rect 193989 149745 209259 149773
rect 209287 149745 209321 149773
rect 209349 149745 224619 149773
rect 224647 149745 224681 149773
rect 224709 149745 239979 149773
rect 240007 149745 240041 149773
rect 240069 149745 256437 149773
rect 256465 149745 256499 149773
rect 256527 149745 256561 149773
rect 256589 149745 256623 149773
rect 256651 149745 265437 149773
rect 265465 149745 265499 149773
rect 265527 149745 265561 149773
rect 265589 149745 265623 149773
rect 265651 149745 274437 149773
rect 274465 149745 274499 149773
rect 274527 149745 274561 149773
rect 274589 149745 274623 149773
rect 274651 149745 283437 149773
rect 283465 149745 283499 149773
rect 283527 149745 283561 149773
rect 283589 149745 283623 149773
rect 283651 149745 292437 149773
rect 292465 149745 292499 149773
rect 292527 149745 292561 149773
rect 292589 149745 292623 149773
rect 292651 149745 299736 149773
rect 299764 149745 299798 149773
rect 299826 149745 299860 149773
rect 299888 149745 299922 149773
rect 299950 149745 299998 149773
rect -6 149697 299998 149745
rect -6 146959 299998 147007
rect -6 146931 522 146959
rect 550 146931 584 146959
rect 612 146931 646 146959
rect 674 146931 708 146959
rect 736 146931 2577 146959
rect 2605 146931 2639 146959
rect 2667 146931 2701 146959
rect 2729 146931 2763 146959
rect 2791 146931 11577 146959
rect 11605 146931 11639 146959
rect 11667 146931 11701 146959
rect 11729 146931 11763 146959
rect 11791 146931 17259 146959
rect 17287 146931 17321 146959
rect 17349 146931 20577 146959
rect 20605 146931 20639 146959
rect 20667 146931 20701 146959
rect 20729 146931 20763 146959
rect 20791 146931 29577 146959
rect 29605 146931 29639 146959
rect 29667 146931 29701 146959
rect 29729 146931 29763 146959
rect 29791 146931 32619 146959
rect 32647 146931 32681 146959
rect 32709 146931 47979 146959
rect 48007 146931 48041 146959
rect 48069 146931 63339 146959
rect 63367 146931 63401 146959
rect 63429 146931 78699 146959
rect 78727 146931 78761 146959
rect 78789 146931 94059 146959
rect 94087 146931 94121 146959
rect 94149 146931 109419 146959
rect 109447 146931 109481 146959
rect 109509 146931 124779 146959
rect 124807 146931 124841 146959
rect 124869 146931 140139 146959
rect 140167 146931 140201 146959
rect 140229 146931 155499 146959
rect 155527 146931 155561 146959
rect 155589 146931 170859 146959
rect 170887 146931 170921 146959
rect 170949 146931 186219 146959
rect 186247 146931 186281 146959
rect 186309 146931 201579 146959
rect 201607 146931 201641 146959
rect 201669 146931 216939 146959
rect 216967 146931 217001 146959
rect 217029 146931 232299 146959
rect 232327 146931 232361 146959
rect 232389 146931 247659 146959
rect 247687 146931 247721 146959
rect 247749 146931 254577 146959
rect 254605 146931 254639 146959
rect 254667 146931 254701 146959
rect 254729 146931 254763 146959
rect 254791 146931 263577 146959
rect 263605 146931 263639 146959
rect 263667 146931 263701 146959
rect 263729 146931 263763 146959
rect 263791 146931 272577 146959
rect 272605 146931 272639 146959
rect 272667 146931 272701 146959
rect 272729 146931 272763 146959
rect 272791 146931 281577 146959
rect 281605 146931 281639 146959
rect 281667 146931 281701 146959
rect 281729 146931 281763 146959
rect 281791 146931 290577 146959
rect 290605 146931 290639 146959
rect 290667 146931 290701 146959
rect 290729 146931 290763 146959
rect 290791 146931 299256 146959
rect 299284 146931 299318 146959
rect 299346 146931 299380 146959
rect 299408 146931 299442 146959
rect 299470 146931 299998 146959
rect -6 146897 299998 146931
rect -6 146869 522 146897
rect 550 146869 584 146897
rect 612 146869 646 146897
rect 674 146869 708 146897
rect 736 146869 2577 146897
rect 2605 146869 2639 146897
rect 2667 146869 2701 146897
rect 2729 146869 2763 146897
rect 2791 146869 11577 146897
rect 11605 146869 11639 146897
rect 11667 146869 11701 146897
rect 11729 146869 11763 146897
rect 11791 146869 17259 146897
rect 17287 146869 17321 146897
rect 17349 146869 20577 146897
rect 20605 146869 20639 146897
rect 20667 146869 20701 146897
rect 20729 146869 20763 146897
rect 20791 146869 29577 146897
rect 29605 146869 29639 146897
rect 29667 146869 29701 146897
rect 29729 146869 29763 146897
rect 29791 146869 32619 146897
rect 32647 146869 32681 146897
rect 32709 146869 47979 146897
rect 48007 146869 48041 146897
rect 48069 146869 63339 146897
rect 63367 146869 63401 146897
rect 63429 146869 78699 146897
rect 78727 146869 78761 146897
rect 78789 146869 94059 146897
rect 94087 146869 94121 146897
rect 94149 146869 109419 146897
rect 109447 146869 109481 146897
rect 109509 146869 124779 146897
rect 124807 146869 124841 146897
rect 124869 146869 140139 146897
rect 140167 146869 140201 146897
rect 140229 146869 155499 146897
rect 155527 146869 155561 146897
rect 155589 146869 170859 146897
rect 170887 146869 170921 146897
rect 170949 146869 186219 146897
rect 186247 146869 186281 146897
rect 186309 146869 201579 146897
rect 201607 146869 201641 146897
rect 201669 146869 216939 146897
rect 216967 146869 217001 146897
rect 217029 146869 232299 146897
rect 232327 146869 232361 146897
rect 232389 146869 247659 146897
rect 247687 146869 247721 146897
rect 247749 146869 254577 146897
rect 254605 146869 254639 146897
rect 254667 146869 254701 146897
rect 254729 146869 254763 146897
rect 254791 146869 263577 146897
rect 263605 146869 263639 146897
rect 263667 146869 263701 146897
rect 263729 146869 263763 146897
rect 263791 146869 272577 146897
rect 272605 146869 272639 146897
rect 272667 146869 272701 146897
rect 272729 146869 272763 146897
rect 272791 146869 281577 146897
rect 281605 146869 281639 146897
rect 281667 146869 281701 146897
rect 281729 146869 281763 146897
rect 281791 146869 290577 146897
rect 290605 146869 290639 146897
rect 290667 146869 290701 146897
rect 290729 146869 290763 146897
rect 290791 146869 299256 146897
rect 299284 146869 299318 146897
rect 299346 146869 299380 146897
rect 299408 146869 299442 146897
rect 299470 146869 299998 146897
rect -6 146835 299998 146869
rect -6 146807 522 146835
rect 550 146807 584 146835
rect 612 146807 646 146835
rect 674 146807 708 146835
rect 736 146807 2577 146835
rect 2605 146807 2639 146835
rect 2667 146807 2701 146835
rect 2729 146807 2763 146835
rect 2791 146807 11577 146835
rect 11605 146807 11639 146835
rect 11667 146807 11701 146835
rect 11729 146807 11763 146835
rect 11791 146807 17259 146835
rect 17287 146807 17321 146835
rect 17349 146807 20577 146835
rect 20605 146807 20639 146835
rect 20667 146807 20701 146835
rect 20729 146807 20763 146835
rect 20791 146807 29577 146835
rect 29605 146807 29639 146835
rect 29667 146807 29701 146835
rect 29729 146807 29763 146835
rect 29791 146807 32619 146835
rect 32647 146807 32681 146835
rect 32709 146807 47979 146835
rect 48007 146807 48041 146835
rect 48069 146807 63339 146835
rect 63367 146807 63401 146835
rect 63429 146807 78699 146835
rect 78727 146807 78761 146835
rect 78789 146807 94059 146835
rect 94087 146807 94121 146835
rect 94149 146807 109419 146835
rect 109447 146807 109481 146835
rect 109509 146807 124779 146835
rect 124807 146807 124841 146835
rect 124869 146807 140139 146835
rect 140167 146807 140201 146835
rect 140229 146807 155499 146835
rect 155527 146807 155561 146835
rect 155589 146807 170859 146835
rect 170887 146807 170921 146835
rect 170949 146807 186219 146835
rect 186247 146807 186281 146835
rect 186309 146807 201579 146835
rect 201607 146807 201641 146835
rect 201669 146807 216939 146835
rect 216967 146807 217001 146835
rect 217029 146807 232299 146835
rect 232327 146807 232361 146835
rect 232389 146807 247659 146835
rect 247687 146807 247721 146835
rect 247749 146807 254577 146835
rect 254605 146807 254639 146835
rect 254667 146807 254701 146835
rect 254729 146807 254763 146835
rect 254791 146807 263577 146835
rect 263605 146807 263639 146835
rect 263667 146807 263701 146835
rect 263729 146807 263763 146835
rect 263791 146807 272577 146835
rect 272605 146807 272639 146835
rect 272667 146807 272701 146835
rect 272729 146807 272763 146835
rect 272791 146807 281577 146835
rect 281605 146807 281639 146835
rect 281667 146807 281701 146835
rect 281729 146807 281763 146835
rect 281791 146807 290577 146835
rect 290605 146807 290639 146835
rect 290667 146807 290701 146835
rect 290729 146807 290763 146835
rect 290791 146807 299256 146835
rect 299284 146807 299318 146835
rect 299346 146807 299380 146835
rect 299408 146807 299442 146835
rect 299470 146807 299998 146835
rect -6 146773 299998 146807
rect -6 146745 522 146773
rect 550 146745 584 146773
rect 612 146745 646 146773
rect 674 146745 708 146773
rect 736 146745 2577 146773
rect 2605 146745 2639 146773
rect 2667 146745 2701 146773
rect 2729 146745 2763 146773
rect 2791 146745 11577 146773
rect 11605 146745 11639 146773
rect 11667 146745 11701 146773
rect 11729 146745 11763 146773
rect 11791 146745 17259 146773
rect 17287 146745 17321 146773
rect 17349 146745 20577 146773
rect 20605 146745 20639 146773
rect 20667 146745 20701 146773
rect 20729 146745 20763 146773
rect 20791 146745 29577 146773
rect 29605 146745 29639 146773
rect 29667 146745 29701 146773
rect 29729 146745 29763 146773
rect 29791 146745 32619 146773
rect 32647 146745 32681 146773
rect 32709 146745 47979 146773
rect 48007 146745 48041 146773
rect 48069 146745 63339 146773
rect 63367 146745 63401 146773
rect 63429 146745 78699 146773
rect 78727 146745 78761 146773
rect 78789 146745 94059 146773
rect 94087 146745 94121 146773
rect 94149 146745 109419 146773
rect 109447 146745 109481 146773
rect 109509 146745 124779 146773
rect 124807 146745 124841 146773
rect 124869 146745 140139 146773
rect 140167 146745 140201 146773
rect 140229 146745 155499 146773
rect 155527 146745 155561 146773
rect 155589 146745 170859 146773
rect 170887 146745 170921 146773
rect 170949 146745 186219 146773
rect 186247 146745 186281 146773
rect 186309 146745 201579 146773
rect 201607 146745 201641 146773
rect 201669 146745 216939 146773
rect 216967 146745 217001 146773
rect 217029 146745 232299 146773
rect 232327 146745 232361 146773
rect 232389 146745 247659 146773
rect 247687 146745 247721 146773
rect 247749 146745 254577 146773
rect 254605 146745 254639 146773
rect 254667 146745 254701 146773
rect 254729 146745 254763 146773
rect 254791 146745 263577 146773
rect 263605 146745 263639 146773
rect 263667 146745 263701 146773
rect 263729 146745 263763 146773
rect 263791 146745 272577 146773
rect 272605 146745 272639 146773
rect 272667 146745 272701 146773
rect 272729 146745 272763 146773
rect 272791 146745 281577 146773
rect 281605 146745 281639 146773
rect 281667 146745 281701 146773
rect 281729 146745 281763 146773
rect 281791 146745 290577 146773
rect 290605 146745 290639 146773
rect 290667 146745 290701 146773
rect 290729 146745 290763 146773
rect 290791 146745 299256 146773
rect 299284 146745 299318 146773
rect 299346 146745 299380 146773
rect 299408 146745 299442 146773
rect 299470 146745 299998 146773
rect -6 146697 299998 146745
rect -6 140959 299998 141007
rect -6 140931 42 140959
rect 70 140931 104 140959
rect 132 140931 166 140959
rect 194 140931 228 140959
rect 256 140931 4437 140959
rect 4465 140931 4499 140959
rect 4527 140931 4561 140959
rect 4589 140931 4623 140959
rect 4651 140931 13437 140959
rect 13465 140931 13499 140959
rect 13527 140931 13561 140959
rect 13589 140931 13623 140959
rect 13651 140931 22437 140959
rect 22465 140931 22499 140959
rect 22527 140931 22561 140959
rect 22589 140931 22623 140959
rect 22651 140931 24939 140959
rect 24967 140931 25001 140959
rect 25029 140931 31437 140959
rect 31465 140931 31499 140959
rect 31527 140931 31561 140959
rect 31589 140931 31623 140959
rect 31651 140931 40299 140959
rect 40327 140931 40361 140959
rect 40389 140931 55659 140959
rect 55687 140931 55721 140959
rect 55749 140931 71019 140959
rect 71047 140931 71081 140959
rect 71109 140931 86379 140959
rect 86407 140931 86441 140959
rect 86469 140931 101739 140959
rect 101767 140931 101801 140959
rect 101829 140931 117099 140959
rect 117127 140931 117161 140959
rect 117189 140931 132459 140959
rect 132487 140931 132521 140959
rect 132549 140931 147819 140959
rect 147847 140931 147881 140959
rect 147909 140931 163179 140959
rect 163207 140931 163241 140959
rect 163269 140931 178539 140959
rect 178567 140931 178601 140959
rect 178629 140931 193899 140959
rect 193927 140931 193961 140959
rect 193989 140931 209259 140959
rect 209287 140931 209321 140959
rect 209349 140931 224619 140959
rect 224647 140931 224681 140959
rect 224709 140931 239979 140959
rect 240007 140931 240041 140959
rect 240069 140931 256437 140959
rect 256465 140931 256499 140959
rect 256527 140931 256561 140959
rect 256589 140931 256623 140959
rect 256651 140931 265437 140959
rect 265465 140931 265499 140959
rect 265527 140931 265561 140959
rect 265589 140931 265623 140959
rect 265651 140931 274437 140959
rect 274465 140931 274499 140959
rect 274527 140931 274561 140959
rect 274589 140931 274623 140959
rect 274651 140931 283437 140959
rect 283465 140931 283499 140959
rect 283527 140931 283561 140959
rect 283589 140931 283623 140959
rect 283651 140931 292437 140959
rect 292465 140931 292499 140959
rect 292527 140931 292561 140959
rect 292589 140931 292623 140959
rect 292651 140931 299736 140959
rect 299764 140931 299798 140959
rect 299826 140931 299860 140959
rect 299888 140931 299922 140959
rect 299950 140931 299998 140959
rect -6 140897 299998 140931
rect -6 140869 42 140897
rect 70 140869 104 140897
rect 132 140869 166 140897
rect 194 140869 228 140897
rect 256 140869 4437 140897
rect 4465 140869 4499 140897
rect 4527 140869 4561 140897
rect 4589 140869 4623 140897
rect 4651 140869 13437 140897
rect 13465 140869 13499 140897
rect 13527 140869 13561 140897
rect 13589 140869 13623 140897
rect 13651 140869 22437 140897
rect 22465 140869 22499 140897
rect 22527 140869 22561 140897
rect 22589 140869 22623 140897
rect 22651 140869 24939 140897
rect 24967 140869 25001 140897
rect 25029 140869 31437 140897
rect 31465 140869 31499 140897
rect 31527 140869 31561 140897
rect 31589 140869 31623 140897
rect 31651 140869 40299 140897
rect 40327 140869 40361 140897
rect 40389 140869 55659 140897
rect 55687 140869 55721 140897
rect 55749 140869 71019 140897
rect 71047 140869 71081 140897
rect 71109 140869 86379 140897
rect 86407 140869 86441 140897
rect 86469 140869 101739 140897
rect 101767 140869 101801 140897
rect 101829 140869 117099 140897
rect 117127 140869 117161 140897
rect 117189 140869 132459 140897
rect 132487 140869 132521 140897
rect 132549 140869 147819 140897
rect 147847 140869 147881 140897
rect 147909 140869 163179 140897
rect 163207 140869 163241 140897
rect 163269 140869 178539 140897
rect 178567 140869 178601 140897
rect 178629 140869 193899 140897
rect 193927 140869 193961 140897
rect 193989 140869 209259 140897
rect 209287 140869 209321 140897
rect 209349 140869 224619 140897
rect 224647 140869 224681 140897
rect 224709 140869 239979 140897
rect 240007 140869 240041 140897
rect 240069 140869 256437 140897
rect 256465 140869 256499 140897
rect 256527 140869 256561 140897
rect 256589 140869 256623 140897
rect 256651 140869 265437 140897
rect 265465 140869 265499 140897
rect 265527 140869 265561 140897
rect 265589 140869 265623 140897
rect 265651 140869 274437 140897
rect 274465 140869 274499 140897
rect 274527 140869 274561 140897
rect 274589 140869 274623 140897
rect 274651 140869 283437 140897
rect 283465 140869 283499 140897
rect 283527 140869 283561 140897
rect 283589 140869 283623 140897
rect 283651 140869 292437 140897
rect 292465 140869 292499 140897
rect 292527 140869 292561 140897
rect 292589 140869 292623 140897
rect 292651 140869 299736 140897
rect 299764 140869 299798 140897
rect 299826 140869 299860 140897
rect 299888 140869 299922 140897
rect 299950 140869 299998 140897
rect -6 140835 299998 140869
rect -6 140807 42 140835
rect 70 140807 104 140835
rect 132 140807 166 140835
rect 194 140807 228 140835
rect 256 140807 4437 140835
rect 4465 140807 4499 140835
rect 4527 140807 4561 140835
rect 4589 140807 4623 140835
rect 4651 140807 13437 140835
rect 13465 140807 13499 140835
rect 13527 140807 13561 140835
rect 13589 140807 13623 140835
rect 13651 140807 22437 140835
rect 22465 140807 22499 140835
rect 22527 140807 22561 140835
rect 22589 140807 22623 140835
rect 22651 140807 24939 140835
rect 24967 140807 25001 140835
rect 25029 140807 31437 140835
rect 31465 140807 31499 140835
rect 31527 140807 31561 140835
rect 31589 140807 31623 140835
rect 31651 140807 40299 140835
rect 40327 140807 40361 140835
rect 40389 140807 55659 140835
rect 55687 140807 55721 140835
rect 55749 140807 71019 140835
rect 71047 140807 71081 140835
rect 71109 140807 86379 140835
rect 86407 140807 86441 140835
rect 86469 140807 101739 140835
rect 101767 140807 101801 140835
rect 101829 140807 117099 140835
rect 117127 140807 117161 140835
rect 117189 140807 132459 140835
rect 132487 140807 132521 140835
rect 132549 140807 147819 140835
rect 147847 140807 147881 140835
rect 147909 140807 163179 140835
rect 163207 140807 163241 140835
rect 163269 140807 178539 140835
rect 178567 140807 178601 140835
rect 178629 140807 193899 140835
rect 193927 140807 193961 140835
rect 193989 140807 209259 140835
rect 209287 140807 209321 140835
rect 209349 140807 224619 140835
rect 224647 140807 224681 140835
rect 224709 140807 239979 140835
rect 240007 140807 240041 140835
rect 240069 140807 256437 140835
rect 256465 140807 256499 140835
rect 256527 140807 256561 140835
rect 256589 140807 256623 140835
rect 256651 140807 265437 140835
rect 265465 140807 265499 140835
rect 265527 140807 265561 140835
rect 265589 140807 265623 140835
rect 265651 140807 274437 140835
rect 274465 140807 274499 140835
rect 274527 140807 274561 140835
rect 274589 140807 274623 140835
rect 274651 140807 283437 140835
rect 283465 140807 283499 140835
rect 283527 140807 283561 140835
rect 283589 140807 283623 140835
rect 283651 140807 292437 140835
rect 292465 140807 292499 140835
rect 292527 140807 292561 140835
rect 292589 140807 292623 140835
rect 292651 140807 299736 140835
rect 299764 140807 299798 140835
rect 299826 140807 299860 140835
rect 299888 140807 299922 140835
rect 299950 140807 299998 140835
rect -6 140773 299998 140807
rect -6 140745 42 140773
rect 70 140745 104 140773
rect 132 140745 166 140773
rect 194 140745 228 140773
rect 256 140745 4437 140773
rect 4465 140745 4499 140773
rect 4527 140745 4561 140773
rect 4589 140745 4623 140773
rect 4651 140745 13437 140773
rect 13465 140745 13499 140773
rect 13527 140745 13561 140773
rect 13589 140745 13623 140773
rect 13651 140745 22437 140773
rect 22465 140745 22499 140773
rect 22527 140745 22561 140773
rect 22589 140745 22623 140773
rect 22651 140745 24939 140773
rect 24967 140745 25001 140773
rect 25029 140745 31437 140773
rect 31465 140745 31499 140773
rect 31527 140745 31561 140773
rect 31589 140745 31623 140773
rect 31651 140745 40299 140773
rect 40327 140745 40361 140773
rect 40389 140745 55659 140773
rect 55687 140745 55721 140773
rect 55749 140745 71019 140773
rect 71047 140745 71081 140773
rect 71109 140745 86379 140773
rect 86407 140745 86441 140773
rect 86469 140745 101739 140773
rect 101767 140745 101801 140773
rect 101829 140745 117099 140773
rect 117127 140745 117161 140773
rect 117189 140745 132459 140773
rect 132487 140745 132521 140773
rect 132549 140745 147819 140773
rect 147847 140745 147881 140773
rect 147909 140745 163179 140773
rect 163207 140745 163241 140773
rect 163269 140745 178539 140773
rect 178567 140745 178601 140773
rect 178629 140745 193899 140773
rect 193927 140745 193961 140773
rect 193989 140745 209259 140773
rect 209287 140745 209321 140773
rect 209349 140745 224619 140773
rect 224647 140745 224681 140773
rect 224709 140745 239979 140773
rect 240007 140745 240041 140773
rect 240069 140745 256437 140773
rect 256465 140745 256499 140773
rect 256527 140745 256561 140773
rect 256589 140745 256623 140773
rect 256651 140745 265437 140773
rect 265465 140745 265499 140773
rect 265527 140745 265561 140773
rect 265589 140745 265623 140773
rect 265651 140745 274437 140773
rect 274465 140745 274499 140773
rect 274527 140745 274561 140773
rect 274589 140745 274623 140773
rect 274651 140745 283437 140773
rect 283465 140745 283499 140773
rect 283527 140745 283561 140773
rect 283589 140745 283623 140773
rect 283651 140745 292437 140773
rect 292465 140745 292499 140773
rect 292527 140745 292561 140773
rect 292589 140745 292623 140773
rect 292651 140745 299736 140773
rect 299764 140745 299798 140773
rect 299826 140745 299860 140773
rect 299888 140745 299922 140773
rect 299950 140745 299998 140773
rect -6 140697 299998 140745
rect -6 137959 299998 138007
rect -6 137931 522 137959
rect 550 137931 584 137959
rect 612 137931 646 137959
rect 674 137931 708 137959
rect 736 137931 2577 137959
rect 2605 137931 2639 137959
rect 2667 137931 2701 137959
rect 2729 137931 2763 137959
rect 2791 137931 11577 137959
rect 11605 137931 11639 137959
rect 11667 137931 11701 137959
rect 11729 137931 11763 137959
rect 11791 137931 17259 137959
rect 17287 137931 17321 137959
rect 17349 137931 20577 137959
rect 20605 137931 20639 137959
rect 20667 137931 20701 137959
rect 20729 137931 20763 137959
rect 20791 137931 29577 137959
rect 29605 137931 29639 137959
rect 29667 137931 29701 137959
rect 29729 137931 29763 137959
rect 29791 137931 32619 137959
rect 32647 137931 32681 137959
rect 32709 137931 47979 137959
rect 48007 137931 48041 137959
rect 48069 137931 63339 137959
rect 63367 137931 63401 137959
rect 63429 137931 78699 137959
rect 78727 137931 78761 137959
rect 78789 137931 94059 137959
rect 94087 137931 94121 137959
rect 94149 137931 109419 137959
rect 109447 137931 109481 137959
rect 109509 137931 124779 137959
rect 124807 137931 124841 137959
rect 124869 137931 140139 137959
rect 140167 137931 140201 137959
rect 140229 137931 155499 137959
rect 155527 137931 155561 137959
rect 155589 137931 170859 137959
rect 170887 137931 170921 137959
rect 170949 137931 186219 137959
rect 186247 137931 186281 137959
rect 186309 137931 201579 137959
rect 201607 137931 201641 137959
rect 201669 137931 216939 137959
rect 216967 137931 217001 137959
rect 217029 137931 232299 137959
rect 232327 137931 232361 137959
rect 232389 137931 247659 137959
rect 247687 137931 247721 137959
rect 247749 137931 254577 137959
rect 254605 137931 254639 137959
rect 254667 137931 254701 137959
rect 254729 137931 254763 137959
rect 254791 137931 263577 137959
rect 263605 137931 263639 137959
rect 263667 137931 263701 137959
rect 263729 137931 263763 137959
rect 263791 137931 272577 137959
rect 272605 137931 272639 137959
rect 272667 137931 272701 137959
rect 272729 137931 272763 137959
rect 272791 137931 281577 137959
rect 281605 137931 281639 137959
rect 281667 137931 281701 137959
rect 281729 137931 281763 137959
rect 281791 137931 290577 137959
rect 290605 137931 290639 137959
rect 290667 137931 290701 137959
rect 290729 137931 290763 137959
rect 290791 137931 299256 137959
rect 299284 137931 299318 137959
rect 299346 137931 299380 137959
rect 299408 137931 299442 137959
rect 299470 137931 299998 137959
rect -6 137897 299998 137931
rect -6 137869 522 137897
rect 550 137869 584 137897
rect 612 137869 646 137897
rect 674 137869 708 137897
rect 736 137869 2577 137897
rect 2605 137869 2639 137897
rect 2667 137869 2701 137897
rect 2729 137869 2763 137897
rect 2791 137869 11577 137897
rect 11605 137869 11639 137897
rect 11667 137869 11701 137897
rect 11729 137869 11763 137897
rect 11791 137869 17259 137897
rect 17287 137869 17321 137897
rect 17349 137869 20577 137897
rect 20605 137869 20639 137897
rect 20667 137869 20701 137897
rect 20729 137869 20763 137897
rect 20791 137869 29577 137897
rect 29605 137869 29639 137897
rect 29667 137869 29701 137897
rect 29729 137869 29763 137897
rect 29791 137869 32619 137897
rect 32647 137869 32681 137897
rect 32709 137869 47979 137897
rect 48007 137869 48041 137897
rect 48069 137869 63339 137897
rect 63367 137869 63401 137897
rect 63429 137869 78699 137897
rect 78727 137869 78761 137897
rect 78789 137869 94059 137897
rect 94087 137869 94121 137897
rect 94149 137869 109419 137897
rect 109447 137869 109481 137897
rect 109509 137869 124779 137897
rect 124807 137869 124841 137897
rect 124869 137869 140139 137897
rect 140167 137869 140201 137897
rect 140229 137869 155499 137897
rect 155527 137869 155561 137897
rect 155589 137869 170859 137897
rect 170887 137869 170921 137897
rect 170949 137869 186219 137897
rect 186247 137869 186281 137897
rect 186309 137869 201579 137897
rect 201607 137869 201641 137897
rect 201669 137869 216939 137897
rect 216967 137869 217001 137897
rect 217029 137869 232299 137897
rect 232327 137869 232361 137897
rect 232389 137869 247659 137897
rect 247687 137869 247721 137897
rect 247749 137869 254577 137897
rect 254605 137869 254639 137897
rect 254667 137869 254701 137897
rect 254729 137869 254763 137897
rect 254791 137869 263577 137897
rect 263605 137869 263639 137897
rect 263667 137869 263701 137897
rect 263729 137869 263763 137897
rect 263791 137869 272577 137897
rect 272605 137869 272639 137897
rect 272667 137869 272701 137897
rect 272729 137869 272763 137897
rect 272791 137869 281577 137897
rect 281605 137869 281639 137897
rect 281667 137869 281701 137897
rect 281729 137869 281763 137897
rect 281791 137869 290577 137897
rect 290605 137869 290639 137897
rect 290667 137869 290701 137897
rect 290729 137869 290763 137897
rect 290791 137869 299256 137897
rect 299284 137869 299318 137897
rect 299346 137869 299380 137897
rect 299408 137869 299442 137897
rect 299470 137869 299998 137897
rect -6 137835 299998 137869
rect -6 137807 522 137835
rect 550 137807 584 137835
rect 612 137807 646 137835
rect 674 137807 708 137835
rect 736 137807 2577 137835
rect 2605 137807 2639 137835
rect 2667 137807 2701 137835
rect 2729 137807 2763 137835
rect 2791 137807 11577 137835
rect 11605 137807 11639 137835
rect 11667 137807 11701 137835
rect 11729 137807 11763 137835
rect 11791 137807 17259 137835
rect 17287 137807 17321 137835
rect 17349 137807 20577 137835
rect 20605 137807 20639 137835
rect 20667 137807 20701 137835
rect 20729 137807 20763 137835
rect 20791 137807 29577 137835
rect 29605 137807 29639 137835
rect 29667 137807 29701 137835
rect 29729 137807 29763 137835
rect 29791 137807 32619 137835
rect 32647 137807 32681 137835
rect 32709 137807 47979 137835
rect 48007 137807 48041 137835
rect 48069 137807 63339 137835
rect 63367 137807 63401 137835
rect 63429 137807 78699 137835
rect 78727 137807 78761 137835
rect 78789 137807 94059 137835
rect 94087 137807 94121 137835
rect 94149 137807 109419 137835
rect 109447 137807 109481 137835
rect 109509 137807 124779 137835
rect 124807 137807 124841 137835
rect 124869 137807 140139 137835
rect 140167 137807 140201 137835
rect 140229 137807 155499 137835
rect 155527 137807 155561 137835
rect 155589 137807 170859 137835
rect 170887 137807 170921 137835
rect 170949 137807 186219 137835
rect 186247 137807 186281 137835
rect 186309 137807 201579 137835
rect 201607 137807 201641 137835
rect 201669 137807 216939 137835
rect 216967 137807 217001 137835
rect 217029 137807 232299 137835
rect 232327 137807 232361 137835
rect 232389 137807 247659 137835
rect 247687 137807 247721 137835
rect 247749 137807 254577 137835
rect 254605 137807 254639 137835
rect 254667 137807 254701 137835
rect 254729 137807 254763 137835
rect 254791 137807 263577 137835
rect 263605 137807 263639 137835
rect 263667 137807 263701 137835
rect 263729 137807 263763 137835
rect 263791 137807 272577 137835
rect 272605 137807 272639 137835
rect 272667 137807 272701 137835
rect 272729 137807 272763 137835
rect 272791 137807 281577 137835
rect 281605 137807 281639 137835
rect 281667 137807 281701 137835
rect 281729 137807 281763 137835
rect 281791 137807 290577 137835
rect 290605 137807 290639 137835
rect 290667 137807 290701 137835
rect 290729 137807 290763 137835
rect 290791 137807 299256 137835
rect 299284 137807 299318 137835
rect 299346 137807 299380 137835
rect 299408 137807 299442 137835
rect 299470 137807 299998 137835
rect -6 137773 299998 137807
rect -6 137745 522 137773
rect 550 137745 584 137773
rect 612 137745 646 137773
rect 674 137745 708 137773
rect 736 137745 2577 137773
rect 2605 137745 2639 137773
rect 2667 137745 2701 137773
rect 2729 137745 2763 137773
rect 2791 137745 11577 137773
rect 11605 137745 11639 137773
rect 11667 137745 11701 137773
rect 11729 137745 11763 137773
rect 11791 137745 17259 137773
rect 17287 137745 17321 137773
rect 17349 137745 20577 137773
rect 20605 137745 20639 137773
rect 20667 137745 20701 137773
rect 20729 137745 20763 137773
rect 20791 137745 29577 137773
rect 29605 137745 29639 137773
rect 29667 137745 29701 137773
rect 29729 137745 29763 137773
rect 29791 137745 32619 137773
rect 32647 137745 32681 137773
rect 32709 137745 47979 137773
rect 48007 137745 48041 137773
rect 48069 137745 63339 137773
rect 63367 137745 63401 137773
rect 63429 137745 78699 137773
rect 78727 137745 78761 137773
rect 78789 137745 94059 137773
rect 94087 137745 94121 137773
rect 94149 137745 109419 137773
rect 109447 137745 109481 137773
rect 109509 137745 124779 137773
rect 124807 137745 124841 137773
rect 124869 137745 140139 137773
rect 140167 137745 140201 137773
rect 140229 137745 155499 137773
rect 155527 137745 155561 137773
rect 155589 137745 170859 137773
rect 170887 137745 170921 137773
rect 170949 137745 186219 137773
rect 186247 137745 186281 137773
rect 186309 137745 201579 137773
rect 201607 137745 201641 137773
rect 201669 137745 216939 137773
rect 216967 137745 217001 137773
rect 217029 137745 232299 137773
rect 232327 137745 232361 137773
rect 232389 137745 247659 137773
rect 247687 137745 247721 137773
rect 247749 137745 254577 137773
rect 254605 137745 254639 137773
rect 254667 137745 254701 137773
rect 254729 137745 254763 137773
rect 254791 137745 263577 137773
rect 263605 137745 263639 137773
rect 263667 137745 263701 137773
rect 263729 137745 263763 137773
rect 263791 137745 272577 137773
rect 272605 137745 272639 137773
rect 272667 137745 272701 137773
rect 272729 137745 272763 137773
rect 272791 137745 281577 137773
rect 281605 137745 281639 137773
rect 281667 137745 281701 137773
rect 281729 137745 281763 137773
rect 281791 137745 290577 137773
rect 290605 137745 290639 137773
rect 290667 137745 290701 137773
rect 290729 137745 290763 137773
rect 290791 137745 299256 137773
rect 299284 137745 299318 137773
rect 299346 137745 299380 137773
rect 299408 137745 299442 137773
rect 299470 137745 299998 137773
rect -6 137697 299998 137745
rect -6 131959 299998 132007
rect -6 131931 42 131959
rect 70 131931 104 131959
rect 132 131931 166 131959
rect 194 131931 228 131959
rect 256 131931 4437 131959
rect 4465 131931 4499 131959
rect 4527 131931 4561 131959
rect 4589 131931 4623 131959
rect 4651 131931 13437 131959
rect 13465 131931 13499 131959
rect 13527 131931 13561 131959
rect 13589 131931 13623 131959
rect 13651 131931 22437 131959
rect 22465 131931 22499 131959
rect 22527 131931 22561 131959
rect 22589 131931 22623 131959
rect 22651 131931 24939 131959
rect 24967 131931 25001 131959
rect 25029 131931 31437 131959
rect 31465 131931 31499 131959
rect 31527 131931 31561 131959
rect 31589 131931 31623 131959
rect 31651 131931 40299 131959
rect 40327 131931 40361 131959
rect 40389 131931 55659 131959
rect 55687 131931 55721 131959
rect 55749 131931 71019 131959
rect 71047 131931 71081 131959
rect 71109 131931 86379 131959
rect 86407 131931 86441 131959
rect 86469 131931 101739 131959
rect 101767 131931 101801 131959
rect 101829 131931 117099 131959
rect 117127 131931 117161 131959
rect 117189 131931 132459 131959
rect 132487 131931 132521 131959
rect 132549 131931 147819 131959
rect 147847 131931 147881 131959
rect 147909 131931 163179 131959
rect 163207 131931 163241 131959
rect 163269 131931 178539 131959
rect 178567 131931 178601 131959
rect 178629 131931 193899 131959
rect 193927 131931 193961 131959
rect 193989 131931 209259 131959
rect 209287 131931 209321 131959
rect 209349 131931 224619 131959
rect 224647 131931 224681 131959
rect 224709 131931 239979 131959
rect 240007 131931 240041 131959
rect 240069 131931 256437 131959
rect 256465 131931 256499 131959
rect 256527 131931 256561 131959
rect 256589 131931 256623 131959
rect 256651 131931 265437 131959
rect 265465 131931 265499 131959
rect 265527 131931 265561 131959
rect 265589 131931 265623 131959
rect 265651 131931 274437 131959
rect 274465 131931 274499 131959
rect 274527 131931 274561 131959
rect 274589 131931 274623 131959
rect 274651 131931 283437 131959
rect 283465 131931 283499 131959
rect 283527 131931 283561 131959
rect 283589 131931 283623 131959
rect 283651 131931 292437 131959
rect 292465 131931 292499 131959
rect 292527 131931 292561 131959
rect 292589 131931 292623 131959
rect 292651 131931 299736 131959
rect 299764 131931 299798 131959
rect 299826 131931 299860 131959
rect 299888 131931 299922 131959
rect 299950 131931 299998 131959
rect -6 131897 299998 131931
rect -6 131869 42 131897
rect 70 131869 104 131897
rect 132 131869 166 131897
rect 194 131869 228 131897
rect 256 131869 4437 131897
rect 4465 131869 4499 131897
rect 4527 131869 4561 131897
rect 4589 131869 4623 131897
rect 4651 131869 13437 131897
rect 13465 131869 13499 131897
rect 13527 131869 13561 131897
rect 13589 131869 13623 131897
rect 13651 131869 22437 131897
rect 22465 131869 22499 131897
rect 22527 131869 22561 131897
rect 22589 131869 22623 131897
rect 22651 131869 24939 131897
rect 24967 131869 25001 131897
rect 25029 131869 31437 131897
rect 31465 131869 31499 131897
rect 31527 131869 31561 131897
rect 31589 131869 31623 131897
rect 31651 131869 40299 131897
rect 40327 131869 40361 131897
rect 40389 131869 55659 131897
rect 55687 131869 55721 131897
rect 55749 131869 71019 131897
rect 71047 131869 71081 131897
rect 71109 131869 86379 131897
rect 86407 131869 86441 131897
rect 86469 131869 101739 131897
rect 101767 131869 101801 131897
rect 101829 131869 117099 131897
rect 117127 131869 117161 131897
rect 117189 131869 132459 131897
rect 132487 131869 132521 131897
rect 132549 131869 147819 131897
rect 147847 131869 147881 131897
rect 147909 131869 163179 131897
rect 163207 131869 163241 131897
rect 163269 131869 178539 131897
rect 178567 131869 178601 131897
rect 178629 131869 193899 131897
rect 193927 131869 193961 131897
rect 193989 131869 209259 131897
rect 209287 131869 209321 131897
rect 209349 131869 224619 131897
rect 224647 131869 224681 131897
rect 224709 131869 239979 131897
rect 240007 131869 240041 131897
rect 240069 131869 256437 131897
rect 256465 131869 256499 131897
rect 256527 131869 256561 131897
rect 256589 131869 256623 131897
rect 256651 131869 265437 131897
rect 265465 131869 265499 131897
rect 265527 131869 265561 131897
rect 265589 131869 265623 131897
rect 265651 131869 274437 131897
rect 274465 131869 274499 131897
rect 274527 131869 274561 131897
rect 274589 131869 274623 131897
rect 274651 131869 283437 131897
rect 283465 131869 283499 131897
rect 283527 131869 283561 131897
rect 283589 131869 283623 131897
rect 283651 131869 292437 131897
rect 292465 131869 292499 131897
rect 292527 131869 292561 131897
rect 292589 131869 292623 131897
rect 292651 131869 299736 131897
rect 299764 131869 299798 131897
rect 299826 131869 299860 131897
rect 299888 131869 299922 131897
rect 299950 131869 299998 131897
rect -6 131835 299998 131869
rect -6 131807 42 131835
rect 70 131807 104 131835
rect 132 131807 166 131835
rect 194 131807 228 131835
rect 256 131807 4437 131835
rect 4465 131807 4499 131835
rect 4527 131807 4561 131835
rect 4589 131807 4623 131835
rect 4651 131807 13437 131835
rect 13465 131807 13499 131835
rect 13527 131807 13561 131835
rect 13589 131807 13623 131835
rect 13651 131807 22437 131835
rect 22465 131807 22499 131835
rect 22527 131807 22561 131835
rect 22589 131807 22623 131835
rect 22651 131807 24939 131835
rect 24967 131807 25001 131835
rect 25029 131807 31437 131835
rect 31465 131807 31499 131835
rect 31527 131807 31561 131835
rect 31589 131807 31623 131835
rect 31651 131807 40299 131835
rect 40327 131807 40361 131835
rect 40389 131807 55659 131835
rect 55687 131807 55721 131835
rect 55749 131807 71019 131835
rect 71047 131807 71081 131835
rect 71109 131807 86379 131835
rect 86407 131807 86441 131835
rect 86469 131807 101739 131835
rect 101767 131807 101801 131835
rect 101829 131807 117099 131835
rect 117127 131807 117161 131835
rect 117189 131807 132459 131835
rect 132487 131807 132521 131835
rect 132549 131807 147819 131835
rect 147847 131807 147881 131835
rect 147909 131807 163179 131835
rect 163207 131807 163241 131835
rect 163269 131807 178539 131835
rect 178567 131807 178601 131835
rect 178629 131807 193899 131835
rect 193927 131807 193961 131835
rect 193989 131807 209259 131835
rect 209287 131807 209321 131835
rect 209349 131807 224619 131835
rect 224647 131807 224681 131835
rect 224709 131807 239979 131835
rect 240007 131807 240041 131835
rect 240069 131807 256437 131835
rect 256465 131807 256499 131835
rect 256527 131807 256561 131835
rect 256589 131807 256623 131835
rect 256651 131807 265437 131835
rect 265465 131807 265499 131835
rect 265527 131807 265561 131835
rect 265589 131807 265623 131835
rect 265651 131807 274437 131835
rect 274465 131807 274499 131835
rect 274527 131807 274561 131835
rect 274589 131807 274623 131835
rect 274651 131807 283437 131835
rect 283465 131807 283499 131835
rect 283527 131807 283561 131835
rect 283589 131807 283623 131835
rect 283651 131807 292437 131835
rect 292465 131807 292499 131835
rect 292527 131807 292561 131835
rect 292589 131807 292623 131835
rect 292651 131807 299736 131835
rect 299764 131807 299798 131835
rect 299826 131807 299860 131835
rect 299888 131807 299922 131835
rect 299950 131807 299998 131835
rect -6 131773 299998 131807
rect -6 131745 42 131773
rect 70 131745 104 131773
rect 132 131745 166 131773
rect 194 131745 228 131773
rect 256 131745 4437 131773
rect 4465 131745 4499 131773
rect 4527 131745 4561 131773
rect 4589 131745 4623 131773
rect 4651 131745 13437 131773
rect 13465 131745 13499 131773
rect 13527 131745 13561 131773
rect 13589 131745 13623 131773
rect 13651 131745 22437 131773
rect 22465 131745 22499 131773
rect 22527 131745 22561 131773
rect 22589 131745 22623 131773
rect 22651 131745 24939 131773
rect 24967 131745 25001 131773
rect 25029 131745 31437 131773
rect 31465 131745 31499 131773
rect 31527 131745 31561 131773
rect 31589 131745 31623 131773
rect 31651 131745 40299 131773
rect 40327 131745 40361 131773
rect 40389 131745 55659 131773
rect 55687 131745 55721 131773
rect 55749 131745 71019 131773
rect 71047 131745 71081 131773
rect 71109 131745 86379 131773
rect 86407 131745 86441 131773
rect 86469 131745 101739 131773
rect 101767 131745 101801 131773
rect 101829 131745 117099 131773
rect 117127 131745 117161 131773
rect 117189 131745 132459 131773
rect 132487 131745 132521 131773
rect 132549 131745 147819 131773
rect 147847 131745 147881 131773
rect 147909 131745 163179 131773
rect 163207 131745 163241 131773
rect 163269 131745 178539 131773
rect 178567 131745 178601 131773
rect 178629 131745 193899 131773
rect 193927 131745 193961 131773
rect 193989 131745 209259 131773
rect 209287 131745 209321 131773
rect 209349 131745 224619 131773
rect 224647 131745 224681 131773
rect 224709 131745 239979 131773
rect 240007 131745 240041 131773
rect 240069 131745 256437 131773
rect 256465 131745 256499 131773
rect 256527 131745 256561 131773
rect 256589 131745 256623 131773
rect 256651 131745 265437 131773
rect 265465 131745 265499 131773
rect 265527 131745 265561 131773
rect 265589 131745 265623 131773
rect 265651 131745 274437 131773
rect 274465 131745 274499 131773
rect 274527 131745 274561 131773
rect 274589 131745 274623 131773
rect 274651 131745 283437 131773
rect 283465 131745 283499 131773
rect 283527 131745 283561 131773
rect 283589 131745 283623 131773
rect 283651 131745 292437 131773
rect 292465 131745 292499 131773
rect 292527 131745 292561 131773
rect 292589 131745 292623 131773
rect 292651 131745 299736 131773
rect 299764 131745 299798 131773
rect 299826 131745 299860 131773
rect 299888 131745 299922 131773
rect 299950 131745 299998 131773
rect -6 131697 299998 131745
rect -6 128959 299998 129007
rect -6 128931 522 128959
rect 550 128931 584 128959
rect 612 128931 646 128959
rect 674 128931 708 128959
rect 736 128931 2577 128959
rect 2605 128931 2639 128959
rect 2667 128931 2701 128959
rect 2729 128931 2763 128959
rect 2791 128931 11577 128959
rect 11605 128931 11639 128959
rect 11667 128931 11701 128959
rect 11729 128931 11763 128959
rect 11791 128931 17259 128959
rect 17287 128931 17321 128959
rect 17349 128931 20577 128959
rect 20605 128931 20639 128959
rect 20667 128931 20701 128959
rect 20729 128931 20763 128959
rect 20791 128931 29577 128959
rect 29605 128931 29639 128959
rect 29667 128931 29701 128959
rect 29729 128931 29763 128959
rect 29791 128931 32619 128959
rect 32647 128931 32681 128959
rect 32709 128931 47979 128959
rect 48007 128931 48041 128959
rect 48069 128931 63339 128959
rect 63367 128931 63401 128959
rect 63429 128931 78699 128959
rect 78727 128931 78761 128959
rect 78789 128931 94059 128959
rect 94087 128931 94121 128959
rect 94149 128931 109419 128959
rect 109447 128931 109481 128959
rect 109509 128931 124779 128959
rect 124807 128931 124841 128959
rect 124869 128931 140139 128959
rect 140167 128931 140201 128959
rect 140229 128931 155499 128959
rect 155527 128931 155561 128959
rect 155589 128931 170859 128959
rect 170887 128931 170921 128959
rect 170949 128931 186219 128959
rect 186247 128931 186281 128959
rect 186309 128931 201579 128959
rect 201607 128931 201641 128959
rect 201669 128931 216939 128959
rect 216967 128931 217001 128959
rect 217029 128931 232299 128959
rect 232327 128931 232361 128959
rect 232389 128931 247659 128959
rect 247687 128931 247721 128959
rect 247749 128931 254577 128959
rect 254605 128931 254639 128959
rect 254667 128931 254701 128959
rect 254729 128931 254763 128959
rect 254791 128931 263577 128959
rect 263605 128931 263639 128959
rect 263667 128931 263701 128959
rect 263729 128931 263763 128959
rect 263791 128931 272577 128959
rect 272605 128931 272639 128959
rect 272667 128931 272701 128959
rect 272729 128931 272763 128959
rect 272791 128931 281577 128959
rect 281605 128931 281639 128959
rect 281667 128931 281701 128959
rect 281729 128931 281763 128959
rect 281791 128931 290577 128959
rect 290605 128931 290639 128959
rect 290667 128931 290701 128959
rect 290729 128931 290763 128959
rect 290791 128931 299256 128959
rect 299284 128931 299318 128959
rect 299346 128931 299380 128959
rect 299408 128931 299442 128959
rect 299470 128931 299998 128959
rect -6 128897 299998 128931
rect -6 128869 522 128897
rect 550 128869 584 128897
rect 612 128869 646 128897
rect 674 128869 708 128897
rect 736 128869 2577 128897
rect 2605 128869 2639 128897
rect 2667 128869 2701 128897
rect 2729 128869 2763 128897
rect 2791 128869 11577 128897
rect 11605 128869 11639 128897
rect 11667 128869 11701 128897
rect 11729 128869 11763 128897
rect 11791 128869 17259 128897
rect 17287 128869 17321 128897
rect 17349 128869 20577 128897
rect 20605 128869 20639 128897
rect 20667 128869 20701 128897
rect 20729 128869 20763 128897
rect 20791 128869 29577 128897
rect 29605 128869 29639 128897
rect 29667 128869 29701 128897
rect 29729 128869 29763 128897
rect 29791 128869 32619 128897
rect 32647 128869 32681 128897
rect 32709 128869 47979 128897
rect 48007 128869 48041 128897
rect 48069 128869 63339 128897
rect 63367 128869 63401 128897
rect 63429 128869 78699 128897
rect 78727 128869 78761 128897
rect 78789 128869 94059 128897
rect 94087 128869 94121 128897
rect 94149 128869 109419 128897
rect 109447 128869 109481 128897
rect 109509 128869 124779 128897
rect 124807 128869 124841 128897
rect 124869 128869 140139 128897
rect 140167 128869 140201 128897
rect 140229 128869 155499 128897
rect 155527 128869 155561 128897
rect 155589 128869 170859 128897
rect 170887 128869 170921 128897
rect 170949 128869 186219 128897
rect 186247 128869 186281 128897
rect 186309 128869 201579 128897
rect 201607 128869 201641 128897
rect 201669 128869 216939 128897
rect 216967 128869 217001 128897
rect 217029 128869 232299 128897
rect 232327 128869 232361 128897
rect 232389 128869 247659 128897
rect 247687 128869 247721 128897
rect 247749 128869 254577 128897
rect 254605 128869 254639 128897
rect 254667 128869 254701 128897
rect 254729 128869 254763 128897
rect 254791 128869 263577 128897
rect 263605 128869 263639 128897
rect 263667 128869 263701 128897
rect 263729 128869 263763 128897
rect 263791 128869 272577 128897
rect 272605 128869 272639 128897
rect 272667 128869 272701 128897
rect 272729 128869 272763 128897
rect 272791 128869 281577 128897
rect 281605 128869 281639 128897
rect 281667 128869 281701 128897
rect 281729 128869 281763 128897
rect 281791 128869 290577 128897
rect 290605 128869 290639 128897
rect 290667 128869 290701 128897
rect 290729 128869 290763 128897
rect 290791 128869 299256 128897
rect 299284 128869 299318 128897
rect 299346 128869 299380 128897
rect 299408 128869 299442 128897
rect 299470 128869 299998 128897
rect -6 128835 299998 128869
rect -6 128807 522 128835
rect 550 128807 584 128835
rect 612 128807 646 128835
rect 674 128807 708 128835
rect 736 128807 2577 128835
rect 2605 128807 2639 128835
rect 2667 128807 2701 128835
rect 2729 128807 2763 128835
rect 2791 128807 11577 128835
rect 11605 128807 11639 128835
rect 11667 128807 11701 128835
rect 11729 128807 11763 128835
rect 11791 128807 17259 128835
rect 17287 128807 17321 128835
rect 17349 128807 20577 128835
rect 20605 128807 20639 128835
rect 20667 128807 20701 128835
rect 20729 128807 20763 128835
rect 20791 128807 29577 128835
rect 29605 128807 29639 128835
rect 29667 128807 29701 128835
rect 29729 128807 29763 128835
rect 29791 128807 32619 128835
rect 32647 128807 32681 128835
rect 32709 128807 47979 128835
rect 48007 128807 48041 128835
rect 48069 128807 63339 128835
rect 63367 128807 63401 128835
rect 63429 128807 78699 128835
rect 78727 128807 78761 128835
rect 78789 128807 94059 128835
rect 94087 128807 94121 128835
rect 94149 128807 109419 128835
rect 109447 128807 109481 128835
rect 109509 128807 124779 128835
rect 124807 128807 124841 128835
rect 124869 128807 140139 128835
rect 140167 128807 140201 128835
rect 140229 128807 155499 128835
rect 155527 128807 155561 128835
rect 155589 128807 170859 128835
rect 170887 128807 170921 128835
rect 170949 128807 186219 128835
rect 186247 128807 186281 128835
rect 186309 128807 201579 128835
rect 201607 128807 201641 128835
rect 201669 128807 216939 128835
rect 216967 128807 217001 128835
rect 217029 128807 232299 128835
rect 232327 128807 232361 128835
rect 232389 128807 247659 128835
rect 247687 128807 247721 128835
rect 247749 128807 254577 128835
rect 254605 128807 254639 128835
rect 254667 128807 254701 128835
rect 254729 128807 254763 128835
rect 254791 128807 263577 128835
rect 263605 128807 263639 128835
rect 263667 128807 263701 128835
rect 263729 128807 263763 128835
rect 263791 128807 272577 128835
rect 272605 128807 272639 128835
rect 272667 128807 272701 128835
rect 272729 128807 272763 128835
rect 272791 128807 281577 128835
rect 281605 128807 281639 128835
rect 281667 128807 281701 128835
rect 281729 128807 281763 128835
rect 281791 128807 290577 128835
rect 290605 128807 290639 128835
rect 290667 128807 290701 128835
rect 290729 128807 290763 128835
rect 290791 128807 299256 128835
rect 299284 128807 299318 128835
rect 299346 128807 299380 128835
rect 299408 128807 299442 128835
rect 299470 128807 299998 128835
rect -6 128773 299998 128807
rect -6 128745 522 128773
rect 550 128745 584 128773
rect 612 128745 646 128773
rect 674 128745 708 128773
rect 736 128745 2577 128773
rect 2605 128745 2639 128773
rect 2667 128745 2701 128773
rect 2729 128745 2763 128773
rect 2791 128745 11577 128773
rect 11605 128745 11639 128773
rect 11667 128745 11701 128773
rect 11729 128745 11763 128773
rect 11791 128745 17259 128773
rect 17287 128745 17321 128773
rect 17349 128745 20577 128773
rect 20605 128745 20639 128773
rect 20667 128745 20701 128773
rect 20729 128745 20763 128773
rect 20791 128745 29577 128773
rect 29605 128745 29639 128773
rect 29667 128745 29701 128773
rect 29729 128745 29763 128773
rect 29791 128745 32619 128773
rect 32647 128745 32681 128773
rect 32709 128745 47979 128773
rect 48007 128745 48041 128773
rect 48069 128745 63339 128773
rect 63367 128745 63401 128773
rect 63429 128745 78699 128773
rect 78727 128745 78761 128773
rect 78789 128745 94059 128773
rect 94087 128745 94121 128773
rect 94149 128745 109419 128773
rect 109447 128745 109481 128773
rect 109509 128745 124779 128773
rect 124807 128745 124841 128773
rect 124869 128745 140139 128773
rect 140167 128745 140201 128773
rect 140229 128745 155499 128773
rect 155527 128745 155561 128773
rect 155589 128745 170859 128773
rect 170887 128745 170921 128773
rect 170949 128745 186219 128773
rect 186247 128745 186281 128773
rect 186309 128745 201579 128773
rect 201607 128745 201641 128773
rect 201669 128745 216939 128773
rect 216967 128745 217001 128773
rect 217029 128745 232299 128773
rect 232327 128745 232361 128773
rect 232389 128745 247659 128773
rect 247687 128745 247721 128773
rect 247749 128745 254577 128773
rect 254605 128745 254639 128773
rect 254667 128745 254701 128773
rect 254729 128745 254763 128773
rect 254791 128745 263577 128773
rect 263605 128745 263639 128773
rect 263667 128745 263701 128773
rect 263729 128745 263763 128773
rect 263791 128745 272577 128773
rect 272605 128745 272639 128773
rect 272667 128745 272701 128773
rect 272729 128745 272763 128773
rect 272791 128745 281577 128773
rect 281605 128745 281639 128773
rect 281667 128745 281701 128773
rect 281729 128745 281763 128773
rect 281791 128745 290577 128773
rect 290605 128745 290639 128773
rect 290667 128745 290701 128773
rect 290729 128745 290763 128773
rect 290791 128745 299256 128773
rect 299284 128745 299318 128773
rect 299346 128745 299380 128773
rect 299408 128745 299442 128773
rect 299470 128745 299998 128773
rect -6 128697 299998 128745
rect -6 122959 299998 123007
rect -6 122931 42 122959
rect 70 122931 104 122959
rect 132 122931 166 122959
rect 194 122931 228 122959
rect 256 122931 4437 122959
rect 4465 122931 4499 122959
rect 4527 122931 4561 122959
rect 4589 122931 4623 122959
rect 4651 122931 13437 122959
rect 13465 122931 13499 122959
rect 13527 122931 13561 122959
rect 13589 122931 13623 122959
rect 13651 122931 22437 122959
rect 22465 122931 22499 122959
rect 22527 122931 22561 122959
rect 22589 122931 22623 122959
rect 22651 122931 24939 122959
rect 24967 122931 25001 122959
rect 25029 122931 31437 122959
rect 31465 122931 31499 122959
rect 31527 122931 31561 122959
rect 31589 122931 31623 122959
rect 31651 122931 40299 122959
rect 40327 122931 40361 122959
rect 40389 122931 55659 122959
rect 55687 122931 55721 122959
rect 55749 122931 71019 122959
rect 71047 122931 71081 122959
rect 71109 122931 86379 122959
rect 86407 122931 86441 122959
rect 86469 122931 101739 122959
rect 101767 122931 101801 122959
rect 101829 122931 117099 122959
rect 117127 122931 117161 122959
rect 117189 122931 132459 122959
rect 132487 122931 132521 122959
rect 132549 122931 147819 122959
rect 147847 122931 147881 122959
rect 147909 122931 163179 122959
rect 163207 122931 163241 122959
rect 163269 122931 178539 122959
rect 178567 122931 178601 122959
rect 178629 122931 193899 122959
rect 193927 122931 193961 122959
rect 193989 122931 209259 122959
rect 209287 122931 209321 122959
rect 209349 122931 224619 122959
rect 224647 122931 224681 122959
rect 224709 122931 239979 122959
rect 240007 122931 240041 122959
rect 240069 122931 256437 122959
rect 256465 122931 256499 122959
rect 256527 122931 256561 122959
rect 256589 122931 256623 122959
rect 256651 122931 265437 122959
rect 265465 122931 265499 122959
rect 265527 122931 265561 122959
rect 265589 122931 265623 122959
rect 265651 122931 274437 122959
rect 274465 122931 274499 122959
rect 274527 122931 274561 122959
rect 274589 122931 274623 122959
rect 274651 122931 283437 122959
rect 283465 122931 283499 122959
rect 283527 122931 283561 122959
rect 283589 122931 283623 122959
rect 283651 122931 292437 122959
rect 292465 122931 292499 122959
rect 292527 122931 292561 122959
rect 292589 122931 292623 122959
rect 292651 122931 299736 122959
rect 299764 122931 299798 122959
rect 299826 122931 299860 122959
rect 299888 122931 299922 122959
rect 299950 122931 299998 122959
rect -6 122897 299998 122931
rect -6 122869 42 122897
rect 70 122869 104 122897
rect 132 122869 166 122897
rect 194 122869 228 122897
rect 256 122869 4437 122897
rect 4465 122869 4499 122897
rect 4527 122869 4561 122897
rect 4589 122869 4623 122897
rect 4651 122869 13437 122897
rect 13465 122869 13499 122897
rect 13527 122869 13561 122897
rect 13589 122869 13623 122897
rect 13651 122869 22437 122897
rect 22465 122869 22499 122897
rect 22527 122869 22561 122897
rect 22589 122869 22623 122897
rect 22651 122869 24939 122897
rect 24967 122869 25001 122897
rect 25029 122869 31437 122897
rect 31465 122869 31499 122897
rect 31527 122869 31561 122897
rect 31589 122869 31623 122897
rect 31651 122869 40299 122897
rect 40327 122869 40361 122897
rect 40389 122869 55659 122897
rect 55687 122869 55721 122897
rect 55749 122869 71019 122897
rect 71047 122869 71081 122897
rect 71109 122869 86379 122897
rect 86407 122869 86441 122897
rect 86469 122869 101739 122897
rect 101767 122869 101801 122897
rect 101829 122869 117099 122897
rect 117127 122869 117161 122897
rect 117189 122869 132459 122897
rect 132487 122869 132521 122897
rect 132549 122869 147819 122897
rect 147847 122869 147881 122897
rect 147909 122869 163179 122897
rect 163207 122869 163241 122897
rect 163269 122869 178539 122897
rect 178567 122869 178601 122897
rect 178629 122869 193899 122897
rect 193927 122869 193961 122897
rect 193989 122869 209259 122897
rect 209287 122869 209321 122897
rect 209349 122869 224619 122897
rect 224647 122869 224681 122897
rect 224709 122869 239979 122897
rect 240007 122869 240041 122897
rect 240069 122869 256437 122897
rect 256465 122869 256499 122897
rect 256527 122869 256561 122897
rect 256589 122869 256623 122897
rect 256651 122869 265437 122897
rect 265465 122869 265499 122897
rect 265527 122869 265561 122897
rect 265589 122869 265623 122897
rect 265651 122869 274437 122897
rect 274465 122869 274499 122897
rect 274527 122869 274561 122897
rect 274589 122869 274623 122897
rect 274651 122869 283437 122897
rect 283465 122869 283499 122897
rect 283527 122869 283561 122897
rect 283589 122869 283623 122897
rect 283651 122869 292437 122897
rect 292465 122869 292499 122897
rect 292527 122869 292561 122897
rect 292589 122869 292623 122897
rect 292651 122869 299736 122897
rect 299764 122869 299798 122897
rect 299826 122869 299860 122897
rect 299888 122869 299922 122897
rect 299950 122869 299998 122897
rect -6 122835 299998 122869
rect -6 122807 42 122835
rect 70 122807 104 122835
rect 132 122807 166 122835
rect 194 122807 228 122835
rect 256 122807 4437 122835
rect 4465 122807 4499 122835
rect 4527 122807 4561 122835
rect 4589 122807 4623 122835
rect 4651 122807 13437 122835
rect 13465 122807 13499 122835
rect 13527 122807 13561 122835
rect 13589 122807 13623 122835
rect 13651 122807 22437 122835
rect 22465 122807 22499 122835
rect 22527 122807 22561 122835
rect 22589 122807 22623 122835
rect 22651 122807 24939 122835
rect 24967 122807 25001 122835
rect 25029 122807 31437 122835
rect 31465 122807 31499 122835
rect 31527 122807 31561 122835
rect 31589 122807 31623 122835
rect 31651 122807 40299 122835
rect 40327 122807 40361 122835
rect 40389 122807 55659 122835
rect 55687 122807 55721 122835
rect 55749 122807 71019 122835
rect 71047 122807 71081 122835
rect 71109 122807 86379 122835
rect 86407 122807 86441 122835
rect 86469 122807 101739 122835
rect 101767 122807 101801 122835
rect 101829 122807 117099 122835
rect 117127 122807 117161 122835
rect 117189 122807 132459 122835
rect 132487 122807 132521 122835
rect 132549 122807 147819 122835
rect 147847 122807 147881 122835
rect 147909 122807 163179 122835
rect 163207 122807 163241 122835
rect 163269 122807 178539 122835
rect 178567 122807 178601 122835
rect 178629 122807 193899 122835
rect 193927 122807 193961 122835
rect 193989 122807 209259 122835
rect 209287 122807 209321 122835
rect 209349 122807 224619 122835
rect 224647 122807 224681 122835
rect 224709 122807 239979 122835
rect 240007 122807 240041 122835
rect 240069 122807 256437 122835
rect 256465 122807 256499 122835
rect 256527 122807 256561 122835
rect 256589 122807 256623 122835
rect 256651 122807 265437 122835
rect 265465 122807 265499 122835
rect 265527 122807 265561 122835
rect 265589 122807 265623 122835
rect 265651 122807 274437 122835
rect 274465 122807 274499 122835
rect 274527 122807 274561 122835
rect 274589 122807 274623 122835
rect 274651 122807 283437 122835
rect 283465 122807 283499 122835
rect 283527 122807 283561 122835
rect 283589 122807 283623 122835
rect 283651 122807 292437 122835
rect 292465 122807 292499 122835
rect 292527 122807 292561 122835
rect 292589 122807 292623 122835
rect 292651 122807 299736 122835
rect 299764 122807 299798 122835
rect 299826 122807 299860 122835
rect 299888 122807 299922 122835
rect 299950 122807 299998 122835
rect -6 122773 299998 122807
rect -6 122745 42 122773
rect 70 122745 104 122773
rect 132 122745 166 122773
rect 194 122745 228 122773
rect 256 122745 4437 122773
rect 4465 122745 4499 122773
rect 4527 122745 4561 122773
rect 4589 122745 4623 122773
rect 4651 122745 13437 122773
rect 13465 122745 13499 122773
rect 13527 122745 13561 122773
rect 13589 122745 13623 122773
rect 13651 122745 22437 122773
rect 22465 122745 22499 122773
rect 22527 122745 22561 122773
rect 22589 122745 22623 122773
rect 22651 122745 24939 122773
rect 24967 122745 25001 122773
rect 25029 122745 31437 122773
rect 31465 122745 31499 122773
rect 31527 122745 31561 122773
rect 31589 122745 31623 122773
rect 31651 122745 40299 122773
rect 40327 122745 40361 122773
rect 40389 122745 55659 122773
rect 55687 122745 55721 122773
rect 55749 122745 71019 122773
rect 71047 122745 71081 122773
rect 71109 122745 86379 122773
rect 86407 122745 86441 122773
rect 86469 122745 101739 122773
rect 101767 122745 101801 122773
rect 101829 122745 117099 122773
rect 117127 122745 117161 122773
rect 117189 122745 132459 122773
rect 132487 122745 132521 122773
rect 132549 122745 147819 122773
rect 147847 122745 147881 122773
rect 147909 122745 163179 122773
rect 163207 122745 163241 122773
rect 163269 122745 178539 122773
rect 178567 122745 178601 122773
rect 178629 122745 193899 122773
rect 193927 122745 193961 122773
rect 193989 122745 209259 122773
rect 209287 122745 209321 122773
rect 209349 122745 224619 122773
rect 224647 122745 224681 122773
rect 224709 122745 239979 122773
rect 240007 122745 240041 122773
rect 240069 122745 256437 122773
rect 256465 122745 256499 122773
rect 256527 122745 256561 122773
rect 256589 122745 256623 122773
rect 256651 122745 265437 122773
rect 265465 122745 265499 122773
rect 265527 122745 265561 122773
rect 265589 122745 265623 122773
rect 265651 122745 274437 122773
rect 274465 122745 274499 122773
rect 274527 122745 274561 122773
rect 274589 122745 274623 122773
rect 274651 122745 283437 122773
rect 283465 122745 283499 122773
rect 283527 122745 283561 122773
rect 283589 122745 283623 122773
rect 283651 122745 292437 122773
rect 292465 122745 292499 122773
rect 292527 122745 292561 122773
rect 292589 122745 292623 122773
rect 292651 122745 299736 122773
rect 299764 122745 299798 122773
rect 299826 122745 299860 122773
rect 299888 122745 299922 122773
rect 299950 122745 299998 122773
rect -6 122697 299998 122745
rect -6 119959 299998 120007
rect -6 119931 522 119959
rect 550 119931 584 119959
rect 612 119931 646 119959
rect 674 119931 708 119959
rect 736 119931 2577 119959
rect 2605 119931 2639 119959
rect 2667 119931 2701 119959
rect 2729 119931 2763 119959
rect 2791 119931 11577 119959
rect 11605 119931 11639 119959
rect 11667 119931 11701 119959
rect 11729 119931 11763 119959
rect 11791 119931 17259 119959
rect 17287 119931 17321 119959
rect 17349 119931 20577 119959
rect 20605 119931 20639 119959
rect 20667 119931 20701 119959
rect 20729 119931 20763 119959
rect 20791 119931 29577 119959
rect 29605 119931 29639 119959
rect 29667 119931 29701 119959
rect 29729 119931 29763 119959
rect 29791 119931 32619 119959
rect 32647 119931 32681 119959
rect 32709 119931 47979 119959
rect 48007 119931 48041 119959
rect 48069 119931 63339 119959
rect 63367 119931 63401 119959
rect 63429 119931 78699 119959
rect 78727 119931 78761 119959
rect 78789 119931 94059 119959
rect 94087 119931 94121 119959
rect 94149 119931 109419 119959
rect 109447 119931 109481 119959
rect 109509 119931 124779 119959
rect 124807 119931 124841 119959
rect 124869 119931 140139 119959
rect 140167 119931 140201 119959
rect 140229 119931 155499 119959
rect 155527 119931 155561 119959
rect 155589 119931 170859 119959
rect 170887 119931 170921 119959
rect 170949 119931 186219 119959
rect 186247 119931 186281 119959
rect 186309 119931 201579 119959
rect 201607 119931 201641 119959
rect 201669 119931 216939 119959
rect 216967 119931 217001 119959
rect 217029 119931 232299 119959
rect 232327 119931 232361 119959
rect 232389 119931 247659 119959
rect 247687 119931 247721 119959
rect 247749 119931 254577 119959
rect 254605 119931 254639 119959
rect 254667 119931 254701 119959
rect 254729 119931 254763 119959
rect 254791 119931 263577 119959
rect 263605 119931 263639 119959
rect 263667 119931 263701 119959
rect 263729 119931 263763 119959
rect 263791 119931 272577 119959
rect 272605 119931 272639 119959
rect 272667 119931 272701 119959
rect 272729 119931 272763 119959
rect 272791 119931 281577 119959
rect 281605 119931 281639 119959
rect 281667 119931 281701 119959
rect 281729 119931 281763 119959
rect 281791 119931 290577 119959
rect 290605 119931 290639 119959
rect 290667 119931 290701 119959
rect 290729 119931 290763 119959
rect 290791 119931 299256 119959
rect 299284 119931 299318 119959
rect 299346 119931 299380 119959
rect 299408 119931 299442 119959
rect 299470 119931 299998 119959
rect -6 119897 299998 119931
rect -6 119869 522 119897
rect 550 119869 584 119897
rect 612 119869 646 119897
rect 674 119869 708 119897
rect 736 119869 2577 119897
rect 2605 119869 2639 119897
rect 2667 119869 2701 119897
rect 2729 119869 2763 119897
rect 2791 119869 11577 119897
rect 11605 119869 11639 119897
rect 11667 119869 11701 119897
rect 11729 119869 11763 119897
rect 11791 119869 17259 119897
rect 17287 119869 17321 119897
rect 17349 119869 20577 119897
rect 20605 119869 20639 119897
rect 20667 119869 20701 119897
rect 20729 119869 20763 119897
rect 20791 119869 29577 119897
rect 29605 119869 29639 119897
rect 29667 119869 29701 119897
rect 29729 119869 29763 119897
rect 29791 119869 32619 119897
rect 32647 119869 32681 119897
rect 32709 119869 47979 119897
rect 48007 119869 48041 119897
rect 48069 119869 63339 119897
rect 63367 119869 63401 119897
rect 63429 119869 78699 119897
rect 78727 119869 78761 119897
rect 78789 119869 94059 119897
rect 94087 119869 94121 119897
rect 94149 119869 109419 119897
rect 109447 119869 109481 119897
rect 109509 119869 124779 119897
rect 124807 119869 124841 119897
rect 124869 119869 140139 119897
rect 140167 119869 140201 119897
rect 140229 119869 155499 119897
rect 155527 119869 155561 119897
rect 155589 119869 170859 119897
rect 170887 119869 170921 119897
rect 170949 119869 186219 119897
rect 186247 119869 186281 119897
rect 186309 119869 201579 119897
rect 201607 119869 201641 119897
rect 201669 119869 216939 119897
rect 216967 119869 217001 119897
rect 217029 119869 232299 119897
rect 232327 119869 232361 119897
rect 232389 119869 247659 119897
rect 247687 119869 247721 119897
rect 247749 119869 254577 119897
rect 254605 119869 254639 119897
rect 254667 119869 254701 119897
rect 254729 119869 254763 119897
rect 254791 119869 263577 119897
rect 263605 119869 263639 119897
rect 263667 119869 263701 119897
rect 263729 119869 263763 119897
rect 263791 119869 272577 119897
rect 272605 119869 272639 119897
rect 272667 119869 272701 119897
rect 272729 119869 272763 119897
rect 272791 119869 281577 119897
rect 281605 119869 281639 119897
rect 281667 119869 281701 119897
rect 281729 119869 281763 119897
rect 281791 119869 290577 119897
rect 290605 119869 290639 119897
rect 290667 119869 290701 119897
rect 290729 119869 290763 119897
rect 290791 119869 299256 119897
rect 299284 119869 299318 119897
rect 299346 119869 299380 119897
rect 299408 119869 299442 119897
rect 299470 119869 299998 119897
rect -6 119835 299998 119869
rect -6 119807 522 119835
rect 550 119807 584 119835
rect 612 119807 646 119835
rect 674 119807 708 119835
rect 736 119807 2577 119835
rect 2605 119807 2639 119835
rect 2667 119807 2701 119835
rect 2729 119807 2763 119835
rect 2791 119807 11577 119835
rect 11605 119807 11639 119835
rect 11667 119807 11701 119835
rect 11729 119807 11763 119835
rect 11791 119807 17259 119835
rect 17287 119807 17321 119835
rect 17349 119807 20577 119835
rect 20605 119807 20639 119835
rect 20667 119807 20701 119835
rect 20729 119807 20763 119835
rect 20791 119807 29577 119835
rect 29605 119807 29639 119835
rect 29667 119807 29701 119835
rect 29729 119807 29763 119835
rect 29791 119807 32619 119835
rect 32647 119807 32681 119835
rect 32709 119807 47979 119835
rect 48007 119807 48041 119835
rect 48069 119807 63339 119835
rect 63367 119807 63401 119835
rect 63429 119807 78699 119835
rect 78727 119807 78761 119835
rect 78789 119807 94059 119835
rect 94087 119807 94121 119835
rect 94149 119807 109419 119835
rect 109447 119807 109481 119835
rect 109509 119807 124779 119835
rect 124807 119807 124841 119835
rect 124869 119807 140139 119835
rect 140167 119807 140201 119835
rect 140229 119807 155499 119835
rect 155527 119807 155561 119835
rect 155589 119807 170859 119835
rect 170887 119807 170921 119835
rect 170949 119807 186219 119835
rect 186247 119807 186281 119835
rect 186309 119807 201579 119835
rect 201607 119807 201641 119835
rect 201669 119807 216939 119835
rect 216967 119807 217001 119835
rect 217029 119807 232299 119835
rect 232327 119807 232361 119835
rect 232389 119807 247659 119835
rect 247687 119807 247721 119835
rect 247749 119807 254577 119835
rect 254605 119807 254639 119835
rect 254667 119807 254701 119835
rect 254729 119807 254763 119835
rect 254791 119807 263577 119835
rect 263605 119807 263639 119835
rect 263667 119807 263701 119835
rect 263729 119807 263763 119835
rect 263791 119807 272577 119835
rect 272605 119807 272639 119835
rect 272667 119807 272701 119835
rect 272729 119807 272763 119835
rect 272791 119807 281577 119835
rect 281605 119807 281639 119835
rect 281667 119807 281701 119835
rect 281729 119807 281763 119835
rect 281791 119807 290577 119835
rect 290605 119807 290639 119835
rect 290667 119807 290701 119835
rect 290729 119807 290763 119835
rect 290791 119807 299256 119835
rect 299284 119807 299318 119835
rect 299346 119807 299380 119835
rect 299408 119807 299442 119835
rect 299470 119807 299998 119835
rect -6 119773 299998 119807
rect -6 119745 522 119773
rect 550 119745 584 119773
rect 612 119745 646 119773
rect 674 119745 708 119773
rect 736 119745 2577 119773
rect 2605 119745 2639 119773
rect 2667 119745 2701 119773
rect 2729 119745 2763 119773
rect 2791 119745 11577 119773
rect 11605 119745 11639 119773
rect 11667 119745 11701 119773
rect 11729 119745 11763 119773
rect 11791 119745 17259 119773
rect 17287 119745 17321 119773
rect 17349 119745 20577 119773
rect 20605 119745 20639 119773
rect 20667 119745 20701 119773
rect 20729 119745 20763 119773
rect 20791 119745 29577 119773
rect 29605 119745 29639 119773
rect 29667 119745 29701 119773
rect 29729 119745 29763 119773
rect 29791 119745 32619 119773
rect 32647 119745 32681 119773
rect 32709 119745 47979 119773
rect 48007 119745 48041 119773
rect 48069 119745 63339 119773
rect 63367 119745 63401 119773
rect 63429 119745 78699 119773
rect 78727 119745 78761 119773
rect 78789 119745 94059 119773
rect 94087 119745 94121 119773
rect 94149 119745 109419 119773
rect 109447 119745 109481 119773
rect 109509 119745 124779 119773
rect 124807 119745 124841 119773
rect 124869 119745 140139 119773
rect 140167 119745 140201 119773
rect 140229 119745 155499 119773
rect 155527 119745 155561 119773
rect 155589 119745 170859 119773
rect 170887 119745 170921 119773
rect 170949 119745 186219 119773
rect 186247 119745 186281 119773
rect 186309 119745 201579 119773
rect 201607 119745 201641 119773
rect 201669 119745 216939 119773
rect 216967 119745 217001 119773
rect 217029 119745 232299 119773
rect 232327 119745 232361 119773
rect 232389 119745 247659 119773
rect 247687 119745 247721 119773
rect 247749 119745 254577 119773
rect 254605 119745 254639 119773
rect 254667 119745 254701 119773
rect 254729 119745 254763 119773
rect 254791 119745 263577 119773
rect 263605 119745 263639 119773
rect 263667 119745 263701 119773
rect 263729 119745 263763 119773
rect 263791 119745 272577 119773
rect 272605 119745 272639 119773
rect 272667 119745 272701 119773
rect 272729 119745 272763 119773
rect 272791 119745 281577 119773
rect 281605 119745 281639 119773
rect 281667 119745 281701 119773
rect 281729 119745 281763 119773
rect 281791 119745 290577 119773
rect 290605 119745 290639 119773
rect 290667 119745 290701 119773
rect 290729 119745 290763 119773
rect 290791 119745 299256 119773
rect 299284 119745 299318 119773
rect 299346 119745 299380 119773
rect 299408 119745 299442 119773
rect 299470 119745 299998 119773
rect -6 119697 299998 119745
rect -6 113959 299998 114007
rect -6 113931 42 113959
rect 70 113931 104 113959
rect 132 113931 166 113959
rect 194 113931 228 113959
rect 256 113931 4437 113959
rect 4465 113931 4499 113959
rect 4527 113931 4561 113959
rect 4589 113931 4623 113959
rect 4651 113931 13437 113959
rect 13465 113931 13499 113959
rect 13527 113931 13561 113959
rect 13589 113931 13623 113959
rect 13651 113931 22437 113959
rect 22465 113931 22499 113959
rect 22527 113931 22561 113959
rect 22589 113931 22623 113959
rect 22651 113931 24939 113959
rect 24967 113931 25001 113959
rect 25029 113931 31437 113959
rect 31465 113931 31499 113959
rect 31527 113931 31561 113959
rect 31589 113931 31623 113959
rect 31651 113931 40299 113959
rect 40327 113931 40361 113959
rect 40389 113931 55659 113959
rect 55687 113931 55721 113959
rect 55749 113931 71019 113959
rect 71047 113931 71081 113959
rect 71109 113931 86379 113959
rect 86407 113931 86441 113959
rect 86469 113931 101739 113959
rect 101767 113931 101801 113959
rect 101829 113931 117099 113959
rect 117127 113931 117161 113959
rect 117189 113931 132459 113959
rect 132487 113931 132521 113959
rect 132549 113931 147819 113959
rect 147847 113931 147881 113959
rect 147909 113931 163179 113959
rect 163207 113931 163241 113959
rect 163269 113931 178539 113959
rect 178567 113931 178601 113959
rect 178629 113931 193899 113959
rect 193927 113931 193961 113959
rect 193989 113931 209259 113959
rect 209287 113931 209321 113959
rect 209349 113931 224619 113959
rect 224647 113931 224681 113959
rect 224709 113931 239979 113959
rect 240007 113931 240041 113959
rect 240069 113931 256437 113959
rect 256465 113931 256499 113959
rect 256527 113931 256561 113959
rect 256589 113931 256623 113959
rect 256651 113931 265437 113959
rect 265465 113931 265499 113959
rect 265527 113931 265561 113959
rect 265589 113931 265623 113959
rect 265651 113931 274437 113959
rect 274465 113931 274499 113959
rect 274527 113931 274561 113959
rect 274589 113931 274623 113959
rect 274651 113931 283437 113959
rect 283465 113931 283499 113959
rect 283527 113931 283561 113959
rect 283589 113931 283623 113959
rect 283651 113931 292437 113959
rect 292465 113931 292499 113959
rect 292527 113931 292561 113959
rect 292589 113931 292623 113959
rect 292651 113931 299736 113959
rect 299764 113931 299798 113959
rect 299826 113931 299860 113959
rect 299888 113931 299922 113959
rect 299950 113931 299998 113959
rect -6 113897 299998 113931
rect -6 113869 42 113897
rect 70 113869 104 113897
rect 132 113869 166 113897
rect 194 113869 228 113897
rect 256 113869 4437 113897
rect 4465 113869 4499 113897
rect 4527 113869 4561 113897
rect 4589 113869 4623 113897
rect 4651 113869 13437 113897
rect 13465 113869 13499 113897
rect 13527 113869 13561 113897
rect 13589 113869 13623 113897
rect 13651 113869 22437 113897
rect 22465 113869 22499 113897
rect 22527 113869 22561 113897
rect 22589 113869 22623 113897
rect 22651 113869 24939 113897
rect 24967 113869 25001 113897
rect 25029 113869 31437 113897
rect 31465 113869 31499 113897
rect 31527 113869 31561 113897
rect 31589 113869 31623 113897
rect 31651 113869 40299 113897
rect 40327 113869 40361 113897
rect 40389 113869 55659 113897
rect 55687 113869 55721 113897
rect 55749 113869 71019 113897
rect 71047 113869 71081 113897
rect 71109 113869 86379 113897
rect 86407 113869 86441 113897
rect 86469 113869 101739 113897
rect 101767 113869 101801 113897
rect 101829 113869 117099 113897
rect 117127 113869 117161 113897
rect 117189 113869 132459 113897
rect 132487 113869 132521 113897
rect 132549 113869 147819 113897
rect 147847 113869 147881 113897
rect 147909 113869 163179 113897
rect 163207 113869 163241 113897
rect 163269 113869 178539 113897
rect 178567 113869 178601 113897
rect 178629 113869 193899 113897
rect 193927 113869 193961 113897
rect 193989 113869 209259 113897
rect 209287 113869 209321 113897
rect 209349 113869 224619 113897
rect 224647 113869 224681 113897
rect 224709 113869 239979 113897
rect 240007 113869 240041 113897
rect 240069 113869 256437 113897
rect 256465 113869 256499 113897
rect 256527 113869 256561 113897
rect 256589 113869 256623 113897
rect 256651 113869 265437 113897
rect 265465 113869 265499 113897
rect 265527 113869 265561 113897
rect 265589 113869 265623 113897
rect 265651 113869 274437 113897
rect 274465 113869 274499 113897
rect 274527 113869 274561 113897
rect 274589 113869 274623 113897
rect 274651 113869 283437 113897
rect 283465 113869 283499 113897
rect 283527 113869 283561 113897
rect 283589 113869 283623 113897
rect 283651 113869 292437 113897
rect 292465 113869 292499 113897
rect 292527 113869 292561 113897
rect 292589 113869 292623 113897
rect 292651 113869 299736 113897
rect 299764 113869 299798 113897
rect 299826 113869 299860 113897
rect 299888 113869 299922 113897
rect 299950 113869 299998 113897
rect -6 113835 299998 113869
rect -6 113807 42 113835
rect 70 113807 104 113835
rect 132 113807 166 113835
rect 194 113807 228 113835
rect 256 113807 4437 113835
rect 4465 113807 4499 113835
rect 4527 113807 4561 113835
rect 4589 113807 4623 113835
rect 4651 113807 13437 113835
rect 13465 113807 13499 113835
rect 13527 113807 13561 113835
rect 13589 113807 13623 113835
rect 13651 113807 22437 113835
rect 22465 113807 22499 113835
rect 22527 113807 22561 113835
rect 22589 113807 22623 113835
rect 22651 113807 24939 113835
rect 24967 113807 25001 113835
rect 25029 113807 31437 113835
rect 31465 113807 31499 113835
rect 31527 113807 31561 113835
rect 31589 113807 31623 113835
rect 31651 113807 40299 113835
rect 40327 113807 40361 113835
rect 40389 113807 55659 113835
rect 55687 113807 55721 113835
rect 55749 113807 71019 113835
rect 71047 113807 71081 113835
rect 71109 113807 86379 113835
rect 86407 113807 86441 113835
rect 86469 113807 101739 113835
rect 101767 113807 101801 113835
rect 101829 113807 117099 113835
rect 117127 113807 117161 113835
rect 117189 113807 132459 113835
rect 132487 113807 132521 113835
rect 132549 113807 147819 113835
rect 147847 113807 147881 113835
rect 147909 113807 163179 113835
rect 163207 113807 163241 113835
rect 163269 113807 178539 113835
rect 178567 113807 178601 113835
rect 178629 113807 193899 113835
rect 193927 113807 193961 113835
rect 193989 113807 209259 113835
rect 209287 113807 209321 113835
rect 209349 113807 224619 113835
rect 224647 113807 224681 113835
rect 224709 113807 239979 113835
rect 240007 113807 240041 113835
rect 240069 113807 256437 113835
rect 256465 113807 256499 113835
rect 256527 113807 256561 113835
rect 256589 113807 256623 113835
rect 256651 113807 265437 113835
rect 265465 113807 265499 113835
rect 265527 113807 265561 113835
rect 265589 113807 265623 113835
rect 265651 113807 274437 113835
rect 274465 113807 274499 113835
rect 274527 113807 274561 113835
rect 274589 113807 274623 113835
rect 274651 113807 283437 113835
rect 283465 113807 283499 113835
rect 283527 113807 283561 113835
rect 283589 113807 283623 113835
rect 283651 113807 292437 113835
rect 292465 113807 292499 113835
rect 292527 113807 292561 113835
rect 292589 113807 292623 113835
rect 292651 113807 299736 113835
rect 299764 113807 299798 113835
rect 299826 113807 299860 113835
rect 299888 113807 299922 113835
rect 299950 113807 299998 113835
rect -6 113773 299998 113807
rect -6 113745 42 113773
rect 70 113745 104 113773
rect 132 113745 166 113773
rect 194 113745 228 113773
rect 256 113745 4437 113773
rect 4465 113745 4499 113773
rect 4527 113745 4561 113773
rect 4589 113745 4623 113773
rect 4651 113745 13437 113773
rect 13465 113745 13499 113773
rect 13527 113745 13561 113773
rect 13589 113745 13623 113773
rect 13651 113745 22437 113773
rect 22465 113745 22499 113773
rect 22527 113745 22561 113773
rect 22589 113745 22623 113773
rect 22651 113745 24939 113773
rect 24967 113745 25001 113773
rect 25029 113745 31437 113773
rect 31465 113745 31499 113773
rect 31527 113745 31561 113773
rect 31589 113745 31623 113773
rect 31651 113745 40299 113773
rect 40327 113745 40361 113773
rect 40389 113745 55659 113773
rect 55687 113745 55721 113773
rect 55749 113745 71019 113773
rect 71047 113745 71081 113773
rect 71109 113745 86379 113773
rect 86407 113745 86441 113773
rect 86469 113745 101739 113773
rect 101767 113745 101801 113773
rect 101829 113745 117099 113773
rect 117127 113745 117161 113773
rect 117189 113745 132459 113773
rect 132487 113745 132521 113773
rect 132549 113745 147819 113773
rect 147847 113745 147881 113773
rect 147909 113745 163179 113773
rect 163207 113745 163241 113773
rect 163269 113745 178539 113773
rect 178567 113745 178601 113773
rect 178629 113745 193899 113773
rect 193927 113745 193961 113773
rect 193989 113745 209259 113773
rect 209287 113745 209321 113773
rect 209349 113745 224619 113773
rect 224647 113745 224681 113773
rect 224709 113745 239979 113773
rect 240007 113745 240041 113773
rect 240069 113745 256437 113773
rect 256465 113745 256499 113773
rect 256527 113745 256561 113773
rect 256589 113745 256623 113773
rect 256651 113745 265437 113773
rect 265465 113745 265499 113773
rect 265527 113745 265561 113773
rect 265589 113745 265623 113773
rect 265651 113745 274437 113773
rect 274465 113745 274499 113773
rect 274527 113745 274561 113773
rect 274589 113745 274623 113773
rect 274651 113745 283437 113773
rect 283465 113745 283499 113773
rect 283527 113745 283561 113773
rect 283589 113745 283623 113773
rect 283651 113745 292437 113773
rect 292465 113745 292499 113773
rect 292527 113745 292561 113773
rect 292589 113745 292623 113773
rect 292651 113745 299736 113773
rect 299764 113745 299798 113773
rect 299826 113745 299860 113773
rect 299888 113745 299922 113773
rect 299950 113745 299998 113773
rect -6 113697 299998 113745
rect -6 110959 299998 111007
rect -6 110931 522 110959
rect 550 110931 584 110959
rect 612 110931 646 110959
rect 674 110931 708 110959
rect 736 110931 2577 110959
rect 2605 110931 2639 110959
rect 2667 110931 2701 110959
rect 2729 110931 2763 110959
rect 2791 110931 11577 110959
rect 11605 110931 11639 110959
rect 11667 110931 11701 110959
rect 11729 110931 11763 110959
rect 11791 110931 17259 110959
rect 17287 110931 17321 110959
rect 17349 110931 20577 110959
rect 20605 110931 20639 110959
rect 20667 110931 20701 110959
rect 20729 110931 20763 110959
rect 20791 110931 29577 110959
rect 29605 110931 29639 110959
rect 29667 110931 29701 110959
rect 29729 110931 29763 110959
rect 29791 110931 32619 110959
rect 32647 110931 32681 110959
rect 32709 110931 47979 110959
rect 48007 110931 48041 110959
rect 48069 110931 63339 110959
rect 63367 110931 63401 110959
rect 63429 110931 78699 110959
rect 78727 110931 78761 110959
rect 78789 110931 94059 110959
rect 94087 110931 94121 110959
rect 94149 110931 109419 110959
rect 109447 110931 109481 110959
rect 109509 110931 124779 110959
rect 124807 110931 124841 110959
rect 124869 110931 140139 110959
rect 140167 110931 140201 110959
rect 140229 110931 155499 110959
rect 155527 110931 155561 110959
rect 155589 110931 170859 110959
rect 170887 110931 170921 110959
rect 170949 110931 186219 110959
rect 186247 110931 186281 110959
rect 186309 110931 201579 110959
rect 201607 110931 201641 110959
rect 201669 110931 216939 110959
rect 216967 110931 217001 110959
rect 217029 110931 232299 110959
rect 232327 110931 232361 110959
rect 232389 110931 247659 110959
rect 247687 110931 247721 110959
rect 247749 110931 254577 110959
rect 254605 110931 254639 110959
rect 254667 110931 254701 110959
rect 254729 110931 254763 110959
rect 254791 110931 263577 110959
rect 263605 110931 263639 110959
rect 263667 110931 263701 110959
rect 263729 110931 263763 110959
rect 263791 110931 272577 110959
rect 272605 110931 272639 110959
rect 272667 110931 272701 110959
rect 272729 110931 272763 110959
rect 272791 110931 281577 110959
rect 281605 110931 281639 110959
rect 281667 110931 281701 110959
rect 281729 110931 281763 110959
rect 281791 110931 290577 110959
rect 290605 110931 290639 110959
rect 290667 110931 290701 110959
rect 290729 110931 290763 110959
rect 290791 110931 299256 110959
rect 299284 110931 299318 110959
rect 299346 110931 299380 110959
rect 299408 110931 299442 110959
rect 299470 110931 299998 110959
rect -6 110897 299998 110931
rect -6 110869 522 110897
rect 550 110869 584 110897
rect 612 110869 646 110897
rect 674 110869 708 110897
rect 736 110869 2577 110897
rect 2605 110869 2639 110897
rect 2667 110869 2701 110897
rect 2729 110869 2763 110897
rect 2791 110869 11577 110897
rect 11605 110869 11639 110897
rect 11667 110869 11701 110897
rect 11729 110869 11763 110897
rect 11791 110869 17259 110897
rect 17287 110869 17321 110897
rect 17349 110869 20577 110897
rect 20605 110869 20639 110897
rect 20667 110869 20701 110897
rect 20729 110869 20763 110897
rect 20791 110869 29577 110897
rect 29605 110869 29639 110897
rect 29667 110869 29701 110897
rect 29729 110869 29763 110897
rect 29791 110869 32619 110897
rect 32647 110869 32681 110897
rect 32709 110869 47979 110897
rect 48007 110869 48041 110897
rect 48069 110869 63339 110897
rect 63367 110869 63401 110897
rect 63429 110869 78699 110897
rect 78727 110869 78761 110897
rect 78789 110869 94059 110897
rect 94087 110869 94121 110897
rect 94149 110869 109419 110897
rect 109447 110869 109481 110897
rect 109509 110869 124779 110897
rect 124807 110869 124841 110897
rect 124869 110869 140139 110897
rect 140167 110869 140201 110897
rect 140229 110869 155499 110897
rect 155527 110869 155561 110897
rect 155589 110869 170859 110897
rect 170887 110869 170921 110897
rect 170949 110869 186219 110897
rect 186247 110869 186281 110897
rect 186309 110869 201579 110897
rect 201607 110869 201641 110897
rect 201669 110869 216939 110897
rect 216967 110869 217001 110897
rect 217029 110869 232299 110897
rect 232327 110869 232361 110897
rect 232389 110869 247659 110897
rect 247687 110869 247721 110897
rect 247749 110869 254577 110897
rect 254605 110869 254639 110897
rect 254667 110869 254701 110897
rect 254729 110869 254763 110897
rect 254791 110869 263577 110897
rect 263605 110869 263639 110897
rect 263667 110869 263701 110897
rect 263729 110869 263763 110897
rect 263791 110869 272577 110897
rect 272605 110869 272639 110897
rect 272667 110869 272701 110897
rect 272729 110869 272763 110897
rect 272791 110869 281577 110897
rect 281605 110869 281639 110897
rect 281667 110869 281701 110897
rect 281729 110869 281763 110897
rect 281791 110869 290577 110897
rect 290605 110869 290639 110897
rect 290667 110869 290701 110897
rect 290729 110869 290763 110897
rect 290791 110869 299256 110897
rect 299284 110869 299318 110897
rect 299346 110869 299380 110897
rect 299408 110869 299442 110897
rect 299470 110869 299998 110897
rect -6 110835 299998 110869
rect -6 110807 522 110835
rect 550 110807 584 110835
rect 612 110807 646 110835
rect 674 110807 708 110835
rect 736 110807 2577 110835
rect 2605 110807 2639 110835
rect 2667 110807 2701 110835
rect 2729 110807 2763 110835
rect 2791 110807 11577 110835
rect 11605 110807 11639 110835
rect 11667 110807 11701 110835
rect 11729 110807 11763 110835
rect 11791 110807 17259 110835
rect 17287 110807 17321 110835
rect 17349 110807 20577 110835
rect 20605 110807 20639 110835
rect 20667 110807 20701 110835
rect 20729 110807 20763 110835
rect 20791 110807 29577 110835
rect 29605 110807 29639 110835
rect 29667 110807 29701 110835
rect 29729 110807 29763 110835
rect 29791 110807 32619 110835
rect 32647 110807 32681 110835
rect 32709 110807 47979 110835
rect 48007 110807 48041 110835
rect 48069 110807 63339 110835
rect 63367 110807 63401 110835
rect 63429 110807 78699 110835
rect 78727 110807 78761 110835
rect 78789 110807 94059 110835
rect 94087 110807 94121 110835
rect 94149 110807 109419 110835
rect 109447 110807 109481 110835
rect 109509 110807 124779 110835
rect 124807 110807 124841 110835
rect 124869 110807 140139 110835
rect 140167 110807 140201 110835
rect 140229 110807 155499 110835
rect 155527 110807 155561 110835
rect 155589 110807 170859 110835
rect 170887 110807 170921 110835
rect 170949 110807 186219 110835
rect 186247 110807 186281 110835
rect 186309 110807 201579 110835
rect 201607 110807 201641 110835
rect 201669 110807 216939 110835
rect 216967 110807 217001 110835
rect 217029 110807 232299 110835
rect 232327 110807 232361 110835
rect 232389 110807 247659 110835
rect 247687 110807 247721 110835
rect 247749 110807 254577 110835
rect 254605 110807 254639 110835
rect 254667 110807 254701 110835
rect 254729 110807 254763 110835
rect 254791 110807 263577 110835
rect 263605 110807 263639 110835
rect 263667 110807 263701 110835
rect 263729 110807 263763 110835
rect 263791 110807 272577 110835
rect 272605 110807 272639 110835
rect 272667 110807 272701 110835
rect 272729 110807 272763 110835
rect 272791 110807 281577 110835
rect 281605 110807 281639 110835
rect 281667 110807 281701 110835
rect 281729 110807 281763 110835
rect 281791 110807 290577 110835
rect 290605 110807 290639 110835
rect 290667 110807 290701 110835
rect 290729 110807 290763 110835
rect 290791 110807 299256 110835
rect 299284 110807 299318 110835
rect 299346 110807 299380 110835
rect 299408 110807 299442 110835
rect 299470 110807 299998 110835
rect -6 110773 299998 110807
rect -6 110745 522 110773
rect 550 110745 584 110773
rect 612 110745 646 110773
rect 674 110745 708 110773
rect 736 110745 2577 110773
rect 2605 110745 2639 110773
rect 2667 110745 2701 110773
rect 2729 110745 2763 110773
rect 2791 110745 11577 110773
rect 11605 110745 11639 110773
rect 11667 110745 11701 110773
rect 11729 110745 11763 110773
rect 11791 110745 17259 110773
rect 17287 110745 17321 110773
rect 17349 110745 20577 110773
rect 20605 110745 20639 110773
rect 20667 110745 20701 110773
rect 20729 110745 20763 110773
rect 20791 110745 29577 110773
rect 29605 110745 29639 110773
rect 29667 110745 29701 110773
rect 29729 110745 29763 110773
rect 29791 110745 32619 110773
rect 32647 110745 32681 110773
rect 32709 110745 47979 110773
rect 48007 110745 48041 110773
rect 48069 110745 63339 110773
rect 63367 110745 63401 110773
rect 63429 110745 78699 110773
rect 78727 110745 78761 110773
rect 78789 110745 94059 110773
rect 94087 110745 94121 110773
rect 94149 110745 109419 110773
rect 109447 110745 109481 110773
rect 109509 110745 124779 110773
rect 124807 110745 124841 110773
rect 124869 110745 140139 110773
rect 140167 110745 140201 110773
rect 140229 110745 155499 110773
rect 155527 110745 155561 110773
rect 155589 110745 170859 110773
rect 170887 110745 170921 110773
rect 170949 110745 186219 110773
rect 186247 110745 186281 110773
rect 186309 110745 201579 110773
rect 201607 110745 201641 110773
rect 201669 110745 216939 110773
rect 216967 110745 217001 110773
rect 217029 110745 232299 110773
rect 232327 110745 232361 110773
rect 232389 110745 247659 110773
rect 247687 110745 247721 110773
rect 247749 110745 254577 110773
rect 254605 110745 254639 110773
rect 254667 110745 254701 110773
rect 254729 110745 254763 110773
rect 254791 110745 263577 110773
rect 263605 110745 263639 110773
rect 263667 110745 263701 110773
rect 263729 110745 263763 110773
rect 263791 110745 272577 110773
rect 272605 110745 272639 110773
rect 272667 110745 272701 110773
rect 272729 110745 272763 110773
rect 272791 110745 281577 110773
rect 281605 110745 281639 110773
rect 281667 110745 281701 110773
rect 281729 110745 281763 110773
rect 281791 110745 290577 110773
rect 290605 110745 290639 110773
rect 290667 110745 290701 110773
rect 290729 110745 290763 110773
rect 290791 110745 299256 110773
rect 299284 110745 299318 110773
rect 299346 110745 299380 110773
rect 299408 110745 299442 110773
rect 299470 110745 299998 110773
rect -6 110697 299998 110745
rect -6 104959 299998 105007
rect -6 104931 42 104959
rect 70 104931 104 104959
rect 132 104931 166 104959
rect 194 104931 228 104959
rect 256 104931 4437 104959
rect 4465 104931 4499 104959
rect 4527 104931 4561 104959
rect 4589 104931 4623 104959
rect 4651 104931 13437 104959
rect 13465 104931 13499 104959
rect 13527 104931 13561 104959
rect 13589 104931 13623 104959
rect 13651 104931 22437 104959
rect 22465 104931 22499 104959
rect 22527 104931 22561 104959
rect 22589 104931 22623 104959
rect 22651 104931 24939 104959
rect 24967 104931 25001 104959
rect 25029 104931 31437 104959
rect 31465 104931 31499 104959
rect 31527 104931 31561 104959
rect 31589 104931 31623 104959
rect 31651 104931 40299 104959
rect 40327 104931 40361 104959
rect 40389 104931 55659 104959
rect 55687 104931 55721 104959
rect 55749 104931 71019 104959
rect 71047 104931 71081 104959
rect 71109 104931 86379 104959
rect 86407 104931 86441 104959
rect 86469 104931 101739 104959
rect 101767 104931 101801 104959
rect 101829 104931 117099 104959
rect 117127 104931 117161 104959
rect 117189 104931 132459 104959
rect 132487 104931 132521 104959
rect 132549 104931 147819 104959
rect 147847 104931 147881 104959
rect 147909 104931 163179 104959
rect 163207 104931 163241 104959
rect 163269 104931 178539 104959
rect 178567 104931 178601 104959
rect 178629 104931 193899 104959
rect 193927 104931 193961 104959
rect 193989 104931 209259 104959
rect 209287 104931 209321 104959
rect 209349 104931 224619 104959
rect 224647 104931 224681 104959
rect 224709 104931 239979 104959
rect 240007 104931 240041 104959
rect 240069 104931 256437 104959
rect 256465 104931 256499 104959
rect 256527 104931 256561 104959
rect 256589 104931 256623 104959
rect 256651 104931 265437 104959
rect 265465 104931 265499 104959
rect 265527 104931 265561 104959
rect 265589 104931 265623 104959
rect 265651 104931 274437 104959
rect 274465 104931 274499 104959
rect 274527 104931 274561 104959
rect 274589 104931 274623 104959
rect 274651 104931 283437 104959
rect 283465 104931 283499 104959
rect 283527 104931 283561 104959
rect 283589 104931 283623 104959
rect 283651 104931 292437 104959
rect 292465 104931 292499 104959
rect 292527 104931 292561 104959
rect 292589 104931 292623 104959
rect 292651 104931 299736 104959
rect 299764 104931 299798 104959
rect 299826 104931 299860 104959
rect 299888 104931 299922 104959
rect 299950 104931 299998 104959
rect -6 104897 299998 104931
rect -6 104869 42 104897
rect 70 104869 104 104897
rect 132 104869 166 104897
rect 194 104869 228 104897
rect 256 104869 4437 104897
rect 4465 104869 4499 104897
rect 4527 104869 4561 104897
rect 4589 104869 4623 104897
rect 4651 104869 13437 104897
rect 13465 104869 13499 104897
rect 13527 104869 13561 104897
rect 13589 104869 13623 104897
rect 13651 104869 22437 104897
rect 22465 104869 22499 104897
rect 22527 104869 22561 104897
rect 22589 104869 22623 104897
rect 22651 104869 24939 104897
rect 24967 104869 25001 104897
rect 25029 104869 31437 104897
rect 31465 104869 31499 104897
rect 31527 104869 31561 104897
rect 31589 104869 31623 104897
rect 31651 104869 40299 104897
rect 40327 104869 40361 104897
rect 40389 104869 55659 104897
rect 55687 104869 55721 104897
rect 55749 104869 71019 104897
rect 71047 104869 71081 104897
rect 71109 104869 86379 104897
rect 86407 104869 86441 104897
rect 86469 104869 101739 104897
rect 101767 104869 101801 104897
rect 101829 104869 117099 104897
rect 117127 104869 117161 104897
rect 117189 104869 132459 104897
rect 132487 104869 132521 104897
rect 132549 104869 147819 104897
rect 147847 104869 147881 104897
rect 147909 104869 163179 104897
rect 163207 104869 163241 104897
rect 163269 104869 178539 104897
rect 178567 104869 178601 104897
rect 178629 104869 193899 104897
rect 193927 104869 193961 104897
rect 193989 104869 209259 104897
rect 209287 104869 209321 104897
rect 209349 104869 224619 104897
rect 224647 104869 224681 104897
rect 224709 104869 239979 104897
rect 240007 104869 240041 104897
rect 240069 104869 256437 104897
rect 256465 104869 256499 104897
rect 256527 104869 256561 104897
rect 256589 104869 256623 104897
rect 256651 104869 265437 104897
rect 265465 104869 265499 104897
rect 265527 104869 265561 104897
rect 265589 104869 265623 104897
rect 265651 104869 274437 104897
rect 274465 104869 274499 104897
rect 274527 104869 274561 104897
rect 274589 104869 274623 104897
rect 274651 104869 283437 104897
rect 283465 104869 283499 104897
rect 283527 104869 283561 104897
rect 283589 104869 283623 104897
rect 283651 104869 292437 104897
rect 292465 104869 292499 104897
rect 292527 104869 292561 104897
rect 292589 104869 292623 104897
rect 292651 104869 299736 104897
rect 299764 104869 299798 104897
rect 299826 104869 299860 104897
rect 299888 104869 299922 104897
rect 299950 104869 299998 104897
rect -6 104835 299998 104869
rect -6 104807 42 104835
rect 70 104807 104 104835
rect 132 104807 166 104835
rect 194 104807 228 104835
rect 256 104807 4437 104835
rect 4465 104807 4499 104835
rect 4527 104807 4561 104835
rect 4589 104807 4623 104835
rect 4651 104807 13437 104835
rect 13465 104807 13499 104835
rect 13527 104807 13561 104835
rect 13589 104807 13623 104835
rect 13651 104807 22437 104835
rect 22465 104807 22499 104835
rect 22527 104807 22561 104835
rect 22589 104807 22623 104835
rect 22651 104807 24939 104835
rect 24967 104807 25001 104835
rect 25029 104807 31437 104835
rect 31465 104807 31499 104835
rect 31527 104807 31561 104835
rect 31589 104807 31623 104835
rect 31651 104807 40299 104835
rect 40327 104807 40361 104835
rect 40389 104807 55659 104835
rect 55687 104807 55721 104835
rect 55749 104807 71019 104835
rect 71047 104807 71081 104835
rect 71109 104807 86379 104835
rect 86407 104807 86441 104835
rect 86469 104807 101739 104835
rect 101767 104807 101801 104835
rect 101829 104807 117099 104835
rect 117127 104807 117161 104835
rect 117189 104807 132459 104835
rect 132487 104807 132521 104835
rect 132549 104807 147819 104835
rect 147847 104807 147881 104835
rect 147909 104807 163179 104835
rect 163207 104807 163241 104835
rect 163269 104807 178539 104835
rect 178567 104807 178601 104835
rect 178629 104807 193899 104835
rect 193927 104807 193961 104835
rect 193989 104807 209259 104835
rect 209287 104807 209321 104835
rect 209349 104807 224619 104835
rect 224647 104807 224681 104835
rect 224709 104807 239979 104835
rect 240007 104807 240041 104835
rect 240069 104807 256437 104835
rect 256465 104807 256499 104835
rect 256527 104807 256561 104835
rect 256589 104807 256623 104835
rect 256651 104807 265437 104835
rect 265465 104807 265499 104835
rect 265527 104807 265561 104835
rect 265589 104807 265623 104835
rect 265651 104807 274437 104835
rect 274465 104807 274499 104835
rect 274527 104807 274561 104835
rect 274589 104807 274623 104835
rect 274651 104807 283437 104835
rect 283465 104807 283499 104835
rect 283527 104807 283561 104835
rect 283589 104807 283623 104835
rect 283651 104807 292437 104835
rect 292465 104807 292499 104835
rect 292527 104807 292561 104835
rect 292589 104807 292623 104835
rect 292651 104807 299736 104835
rect 299764 104807 299798 104835
rect 299826 104807 299860 104835
rect 299888 104807 299922 104835
rect 299950 104807 299998 104835
rect -6 104773 299998 104807
rect -6 104745 42 104773
rect 70 104745 104 104773
rect 132 104745 166 104773
rect 194 104745 228 104773
rect 256 104745 4437 104773
rect 4465 104745 4499 104773
rect 4527 104745 4561 104773
rect 4589 104745 4623 104773
rect 4651 104745 13437 104773
rect 13465 104745 13499 104773
rect 13527 104745 13561 104773
rect 13589 104745 13623 104773
rect 13651 104745 22437 104773
rect 22465 104745 22499 104773
rect 22527 104745 22561 104773
rect 22589 104745 22623 104773
rect 22651 104745 24939 104773
rect 24967 104745 25001 104773
rect 25029 104745 31437 104773
rect 31465 104745 31499 104773
rect 31527 104745 31561 104773
rect 31589 104745 31623 104773
rect 31651 104745 40299 104773
rect 40327 104745 40361 104773
rect 40389 104745 55659 104773
rect 55687 104745 55721 104773
rect 55749 104745 71019 104773
rect 71047 104745 71081 104773
rect 71109 104745 86379 104773
rect 86407 104745 86441 104773
rect 86469 104745 101739 104773
rect 101767 104745 101801 104773
rect 101829 104745 117099 104773
rect 117127 104745 117161 104773
rect 117189 104745 132459 104773
rect 132487 104745 132521 104773
rect 132549 104745 147819 104773
rect 147847 104745 147881 104773
rect 147909 104745 163179 104773
rect 163207 104745 163241 104773
rect 163269 104745 178539 104773
rect 178567 104745 178601 104773
rect 178629 104745 193899 104773
rect 193927 104745 193961 104773
rect 193989 104745 209259 104773
rect 209287 104745 209321 104773
rect 209349 104745 224619 104773
rect 224647 104745 224681 104773
rect 224709 104745 239979 104773
rect 240007 104745 240041 104773
rect 240069 104745 256437 104773
rect 256465 104745 256499 104773
rect 256527 104745 256561 104773
rect 256589 104745 256623 104773
rect 256651 104745 265437 104773
rect 265465 104745 265499 104773
rect 265527 104745 265561 104773
rect 265589 104745 265623 104773
rect 265651 104745 274437 104773
rect 274465 104745 274499 104773
rect 274527 104745 274561 104773
rect 274589 104745 274623 104773
rect 274651 104745 283437 104773
rect 283465 104745 283499 104773
rect 283527 104745 283561 104773
rect 283589 104745 283623 104773
rect 283651 104745 292437 104773
rect 292465 104745 292499 104773
rect 292527 104745 292561 104773
rect 292589 104745 292623 104773
rect 292651 104745 299736 104773
rect 299764 104745 299798 104773
rect 299826 104745 299860 104773
rect 299888 104745 299922 104773
rect 299950 104745 299998 104773
rect -6 104697 299998 104745
rect -6 101959 299998 102007
rect -6 101931 522 101959
rect 550 101931 584 101959
rect 612 101931 646 101959
rect 674 101931 708 101959
rect 736 101931 2577 101959
rect 2605 101931 2639 101959
rect 2667 101931 2701 101959
rect 2729 101931 2763 101959
rect 2791 101931 11577 101959
rect 11605 101931 11639 101959
rect 11667 101931 11701 101959
rect 11729 101931 11763 101959
rect 11791 101931 17259 101959
rect 17287 101931 17321 101959
rect 17349 101931 20577 101959
rect 20605 101931 20639 101959
rect 20667 101931 20701 101959
rect 20729 101931 20763 101959
rect 20791 101931 29577 101959
rect 29605 101931 29639 101959
rect 29667 101931 29701 101959
rect 29729 101931 29763 101959
rect 29791 101931 32619 101959
rect 32647 101931 32681 101959
rect 32709 101931 47979 101959
rect 48007 101931 48041 101959
rect 48069 101931 63339 101959
rect 63367 101931 63401 101959
rect 63429 101931 78699 101959
rect 78727 101931 78761 101959
rect 78789 101931 94059 101959
rect 94087 101931 94121 101959
rect 94149 101931 109419 101959
rect 109447 101931 109481 101959
rect 109509 101931 124779 101959
rect 124807 101931 124841 101959
rect 124869 101931 140139 101959
rect 140167 101931 140201 101959
rect 140229 101931 155499 101959
rect 155527 101931 155561 101959
rect 155589 101931 170859 101959
rect 170887 101931 170921 101959
rect 170949 101931 186219 101959
rect 186247 101931 186281 101959
rect 186309 101931 201579 101959
rect 201607 101931 201641 101959
rect 201669 101931 216939 101959
rect 216967 101931 217001 101959
rect 217029 101931 232299 101959
rect 232327 101931 232361 101959
rect 232389 101931 247659 101959
rect 247687 101931 247721 101959
rect 247749 101931 254577 101959
rect 254605 101931 254639 101959
rect 254667 101931 254701 101959
rect 254729 101931 254763 101959
rect 254791 101931 263577 101959
rect 263605 101931 263639 101959
rect 263667 101931 263701 101959
rect 263729 101931 263763 101959
rect 263791 101931 272577 101959
rect 272605 101931 272639 101959
rect 272667 101931 272701 101959
rect 272729 101931 272763 101959
rect 272791 101931 281577 101959
rect 281605 101931 281639 101959
rect 281667 101931 281701 101959
rect 281729 101931 281763 101959
rect 281791 101931 290577 101959
rect 290605 101931 290639 101959
rect 290667 101931 290701 101959
rect 290729 101931 290763 101959
rect 290791 101931 299256 101959
rect 299284 101931 299318 101959
rect 299346 101931 299380 101959
rect 299408 101931 299442 101959
rect 299470 101931 299998 101959
rect -6 101897 299998 101931
rect -6 101869 522 101897
rect 550 101869 584 101897
rect 612 101869 646 101897
rect 674 101869 708 101897
rect 736 101869 2577 101897
rect 2605 101869 2639 101897
rect 2667 101869 2701 101897
rect 2729 101869 2763 101897
rect 2791 101869 11577 101897
rect 11605 101869 11639 101897
rect 11667 101869 11701 101897
rect 11729 101869 11763 101897
rect 11791 101869 17259 101897
rect 17287 101869 17321 101897
rect 17349 101869 20577 101897
rect 20605 101869 20639 101897
rect 20667 101869 20701 101897
rect 20729 101869 20763 101897
rect 20791 101869 29577 101897
rect 29605 101869 29639 101897
rect 29667 101869 29701 101897
rect 29729 101869 29763 101897
rect 29791 101869 32619 101897
rect 32647 101869 32681 101897
rect 32709 101869 47979 101897
rect 48007 101869 48041 101897
rect 48069 101869 63339 101897
rect 63367 101869 63401 101897
rect 63429 101869 78699 101897
rect 78727 101869 78761 101897
rect 78789 101869 94059 101897
rect 94087 101869 94121 101897
rect 94149 101869 109419 101897
rect 109447 101869 109481 101897
rect 109509 101869 124779 101897
rect 124807 101869 124841 101897
rect 124869 101869 140139 101897
rect 140167 101869 140201 101897
rect 140229 101869 155499 101897
rect 155527 101869 155561 101897
rect 155589 101869 170859 101897
rect 170887 101869 170921 101897
rect 170949 101869 186219 101897
rect 186247 101869 186281 101897
rect 186309 101869 201579 101897
rect 201607 101869 201641 101897
rect 201669 101869 216939 101897
rect 216967 101869 217001 101897
rect 217029 101869 232299 101897
rect 232327 101869 232361 101897
rect 232389 101869 247659 101897
rect 247687 101869 247721 101897
rect 247749 101869 254577 101897
rect 254605 101869 254639 101897
rect 254667 101869 254701 101897
rect 254729 101869 254763 101897
rect 254791 101869 263577 101897
rect 263605 101869 263639 101897
rect 263667 101869 263701 101897
rect 263729 101869 263763 101897
rect 263791 101869 272577 101897
rect 272605 101869 272639 101897
rect 272667 101869 272701 101897
rect 272729 101869 272763 101897
rect 272791 101869 281577 101897
rect 281605 101869 281639 101897
rect 281667 101869 281701 101897
rect 281729 101869 281763 101897
rect 281791 101869 290577 101897
rect 290605 101869 290639 101897
rect 290667 101869 290701 101897
rect 290729 101869 290763 101897
rect 290791 101869 299256 101897
rect 299284 101869 299318 101897
rect 299346 101869 299380 101897
rect 299408 101869 299442 101897
rect 299470 101869 299998 101897
rect -6 101835 299998 101869
rect -6 101807 522 101835
rect 550 101807 584 101835
rect 612 101807 646 101835
rect 674 101807 708 101835
rect 736 101807 2577 101835
rect 2605 101807 2639 101835
rect 2667 101807 2701 101835
rect 2729 101807 2763 101835
rect 2791 101807 11577 101835
rect 11605 101807 11639 101835
rect 11667 101807 11701 101835
rect 11729 101807 11763 101835
rect 11791 101807 17259 101835
rect 17287 101807 17321 101835
rect 17349 101807 20577 101835
rect 20605 101807 20639 101835
rect 20667 101807 20701 101835
rect 20729 101807 20763 101835
rect 20791 101807 29577 101835
rect 29605 101807 29639 101835
rect 29667 101807 29701 101835
rect 29729 101807 29763 101835
rect 29791 101807 32619 101835
rect 32647 101807 32681 101835
rect 32709 101807 47979 101835
rect 48007 101807 48041 101835
rect 48069 101807 63339 101835
rect 63367 101807 63401 101835
rect 63429 101807 78699 101835
rect 78727 101807 78761 101835
rect 78789 101807 94059 101835
rect 94087 101807 94121 101835
rect 94149 101807 109419 101835
rect 109447 101807 109481 101835
rect 109509 101807 124779 101835
rect 124807 101807 124841 101835
rect 124869 101807 140139 101835
rect 140167 101807 140201 101835
rect 140229 101807 155499 101835
rect 155527 101807 155561 101835
rect 155589 101807 170859 101835
rect 170887 101807 170921 101835
rect 170949 101807 186219 101835
rect 186247 101807 186281 101835
rect 186309 101807 201579 101835
rect 201607 101807 201641 101835
rect 201669 101807 216939 101835
rect 216967 101807 217001 101835
rect 217029 101807 232299 101835
rect 232327 101807 232361 101835
rect 232389 101807 247659 101835
rect 247687 101807 247721 101835
rect 247749 101807 254577 101835
rect 254605 101807 254639 101835
rect 254667 101807 254701 101835
rect 254729 101807 254763 101835
rect 254791 101807 263577 101835
rect 263605 101807 263639 101835
rect 263667 101807 263701 101835
rect 263729 101807 263763 101835
rect 263791 101807 272577 101835
rect 272605 101807 272639 101835
rect 272667 101807 272701 101835
rect 272729 101807 272763 101835
rect 272791 101807 281577 101835
rect 281605 101807 281639 101835
rect 281667 101807 281701 101835
rect 281729 101807 281763 101835
rect 281791 101807 290577 101835
rect 290605 101807 290639 101835
rect 290667 101807 290701 101835
rect 290729 101807 290763 101835
rect 290791 101807 299256 101835
rect 299284 101807 299318 101835
rect 299346 101807 299380 101835
rect 299408 101807 299442 101835
rect 299470 101807 299998 101835
rect -6 101773 299998 101807
rect -6 101745 522 101773
rect 550 101745 584 101773
rect 612 101745 646 101773
rect 674 101745 708 101773
rect 736 101745 2577 101773
rect 2605 101745 2639 101773
rect 2667 101745 2701 101773
rect 2729 101745 2763 101773
rect 2791 101745 11577 101773
rect 11605 101745 11639 101773
rect 11667 101745 11701 101773
rect 11729 101745 11763 101773
rect 11791 101745 17259 101773
rect 17287 101745 17321 101773
rect 17349 101745 20577 101773
rect 20605 101745 20639 101773
rect 20667 101745 20701 101773
rect 20729 101745 20763 101773
rect 20791 101745 29577 101773
rect 29605 101745 29639 101773
rect 29667 101745 29701 101773
rect 29729 101745 29763 101773
rect 29791 101745 32619 101773
rect 32647 101745 32681 101773
rect 32709 101745 47979 101773
rect 48007 101745 48041 101773
rect 48069 101745 63339 101773
rect 63367 101745 63401 101773
rect 63429 101745 78699 101773
rect 78727 101745 78761 101773
rect 78789 101745 94059 101773
rect 94087 101745 94121 101773
rect 94149 101745 109419 101773
rect 109447 101745 109481 101773
rect 109509 101745 124779 101773
rect 124807 101745 124841 101773
rect 124869 101745 140139 101773
rect 140167 101745 140201 101773
rect 140229 101745 155499 101773
rect 155527 101745 155561 101773
rect 155589 101745 170859 101773
rect 170887 101745 170921 101773
rect 170949 101745 186219 101773
rect 186247 101745 186281 101773
rect 186309 101745 201579 101773
rect 201607 101745 201641 101773
rect 201669 101745 216939 101773
rect 216967 101745 217001 101773
rect 217029 101745 232299 101773
rect 232327 101745 232361 101773
rect 232389 101745 247659 101773
rect 247687 101745 247721 101773
rect 247749 101745 254577 101773
rect 254605 101745 254639 101773
rect 254667 101745 254701 101773
rect 254729 101745 254763 101773
rect 254791 101745 263577 101773
rect 263605 101745 263639 101773
rect 263667 101745 263701 101773
rect 263729 101745 263763 101773
rect 263791 101745 272577 101773
rect 272605 101745 272639 101773
rect 272667 101745 272701 101773
rect 272729 101745 272763 101773
rect 272791 101745 281577 101773
rect 281605 101745 281639 101773
rect 281667 101745 281701 101773
rect 281729 101745 281763 101773
rect 281791 101745 290577 101773
rect 290605 101745 290639 101773
rect 290667 101745 290701 101773
rect 290729 101745 290763 101773
rect 290791 101745 299256 101773
rect 299284 101745 299318 101773
rect 299346 101745 299380 101773
rect 299408 101745 299442 101773
rect 299470 101745 299998 101773
rect -6 101697 299998 101745
rect -6 95959 299998 96007
rect -6 95931 42 95959
rect 70 95931 104 95959
rect 132 95931 166 95959
rect 194 95931 228 95959
rect 256 95931 4437 95959
rect 4465 95931 4499 95959
rect 4527 95931 4561 95959
rect 4589 95931 4623 95959
rect 4651 95931 13437 95959
rect 13465 95931 13499 95959
rect 13527 95931 13561 95959
rect 13589 95931 13623 95959
rect 13651 95931 22437 95959
rect 22465 95931 22499 95959
rect 22527 95931 22561 95959
rect 22589 95931 22623 95959
rect 22651 95931 24939 95959
rect 24967 95931 25001 95959
rect 25029 95931 31437 95959
rect 31465 95931 31499 95959
rect 31527 95931 31561 95959
rect 31589 95931 31623 95959
rect 31651 95931 40299 95959
rect 40327 95931 40361 95959
rect 40389 95931 55659 95959
rect 55687 95931 55721 95959
rect 55749 95931 71019 95959
rect 71047 95931 71081 95959
rect 71109 95931 86379 95959
rect 86407 95931 86441 95959
rect 86469 95931 101739 95959
rect 101767 95931 101801 95959
rect 101829 95931 117099 95959
rect 117127 95931 117161 95959
rect 117189 95931 132459 95959
rect 132487 95931 132521 95959
rect 132549 95931 147819 95959
rect 147847 95931 147881 95959
rect 147909 95931 163179 95959
rect 163207 95931 163241 95959
rect 163269 95931 178539 95959
rect 178567 95931 178601 95959
rect 178629 95931 193899 95959
rect 193927 95931 193961 95959
rect 193989 95931 209259 95959
rect 209287 95931 209321 95959
rect 209349 95931 224619 95959
rect 224647 95931 224681 95959
rect 224709 95931 239979 95959
rect 240007 95931 240041 95959
rect 240069 95931 256437 95959
rect 256465 95931 256499 95959
rect 256527 95931 256561 95959
rect 256589 95931 256623 95959
rect 256651 95931 265437 95959
rect 265465 95931 265499 95959
rect 265527 95931 265561 95959
rect 265589 95931 265623 95959
rect 265651 95931 274437 95959
rect 274465 95931 274499 95959
rect 274527 95931 274561 95959
rect 274589 95931 274623 95959
rect 274651 95931 283437 95959
rect 283465 95931 283499 95959
rect 283527 95931 283561 95959
rect 283589 95931 283623 95959
rect 283651 95931 292437 95959
rect 292465 95931 292499 95959
rect 292527 95931 292561 95959
rect 292589 95931 292623 95959
rect 292651 95931 299736 95959
rect 299764 95931 299798 95959
rect 299826 95931 299860 95959
rect 299888 95931 299922 95959
rect 299950 95931 299998 95959
rect -6 95897 299998 95931
rect -6 95869 42 95897
rect 70 95869 104 95897
rect 132 95869 166 95897
rect 194 95869 228 95897
rect 256 95869 4437 95897
rect 4465 95869 4499 95897
rect 4527 95869 4561 95897
rect 4589 95869 4623 95897
rect 4651 95869 13437 95897
rect 13465 95869 13499 95897
rect 13527 95869 13561 95897
rect 13589 95869 13623 95897
rect 13651 95869 22437 95897
rect 22465 95869 22499 95897
rect 22527 95869 22561 95897
rect 22589 95869 22623 95897
rect 22651 95869 24939 95897
rect 24967 95869 25001 95897
rect 25029 95869 31437 95897
rect 31465 95869 31499 95897
rect 31527 95869 31561 95897
rect 31589 95869 31623 95897
rect 31651 95869 40299 95897
rect 40327 95869 40361 95897
rect 40389 95869 55659 95897
rect 55687 95869 55721 95897
rect 55749 95869 71019 95897
rect 71047 95869 71081 95897
rect 71109 95869 86379 95897
rect 86407 95869 86441 95897
rect 86469 95869 101739 95897
rect 101767 95869 101801 95897
rect 101829 95869 117099 95897
rect 117127 95869 117161 95897
rect 117189 95869 132459 95897
rect 132487 95869 132521 95897
rect 132549 95869 147819 95897
rect 147847 95869 147881 95897
rect 147909 95869 163179 95897
rect 163207 95869 163241 95897
rect 163269 95869 178539 95897
rect 178567 95869 178601 95897
rect 178629 95869 193899 95897
rect 193927 95869 193961 95897
rect 193989 95869 209259 95897
rect 209287 95869 209321 95897
rect 209349 95869 224619 95897
rect 224647 95869 224681 95897
rect 224709 95869 239979 95897
rect 240007 95869 240041 95897
rect 240069 95869 256437 95897
rect 256465 95869 256499 95897
rect 256527 95869 256561 95897
rect 256589 95869 256623 95897
rect 256651 95869 265437 95897
rect 265465 95869 265499 95897
rect 265527 95869 265561 95897
rect 265589 95869 265623 95897
rect 265651 95869 274437 95897
rect 274465 95869 274499 95897
rect 274527 95869 274561 95897
rect 274589 95869 274623 95897
rect 274651 95869 283437 95897
rect 283465 95869 283499 95897
rect 283527 95869 283561 95897
rect 283589 95869 283623 95897
rect 283651 95869 292437 95897
rect 292465 95869 292499 95897
rect 292527 95869 292561 95897
rect 292589 95869 292623 95897
rect 292651 95869 299736 95897
rect 299764 95869 299798 95897
rect 299826 95869 299860 95897
rect 299888 95869 299922 95897
rect 299950 95869 299998 95897
rect -6 95835 299998 95869
rect -6 95807 42 95835
rect 70 95807 104 95835
rect 132 95807 166 95835
rect 194 95807 228 95835
rect 256 95807 4437 95835
rect 4465 95807 4499 95835
rect 4527 95807 4561 95835
rect 4589 95807 4623 95835
rect 4651 95807 13437 95835
rect 13465 95807 13499 95835
rect 13527 95807 13561 95835
rect 13589 95807 13623 95835
rect 13651 95807 22437 95835
rect 22465 95807 22499 95835
rect 22527 95807 22561 95835
rect 22589 95807 22623 95835
rect 22651 95807 24939 95835
rect 24967 95807 25001 95835
rect 25029 95807 31437 95835
rect 31465 95807 31499 95835
rect 31527 95807 31561 95835
rect 31589 95807 31623 95835
rect 31651 95807 40299 95835
rect 40327 95807 40361 95835
rect 40389 95807 55659 95835
rect 55687 95807 55721 95835
rect 55749 95807 71019 95835
rect 71047 95807 71081 95835
rect 71109 95807 86379 95835
rect 86407 95807 86441 95835
rect 86469 95807 101739 95835
rect 101767 95807 101801 95835
rect 101829 95807 117099 95835
rect 117127 95807 117161 95835
rect 117189 95807 132459 95835
rect 132487 95807 132521 95835
rect 132549 95807 147819 95835
rect 147847 95807 147881 95835
rect 147909 95807 163179 95835
rect 163207 95807 163241 95835
rect 163269 95807 178539 95835
rect 178567 95807 178601 95835
rect 178629 95807 193899 95835
rect 193927 95807 193961 95835
rect 193989 95807 209259 95835
rect 209287 95807 209321 95835
rect 209349 95807 224619 95835
rect 224647 95807 224681 95835
rect 224709 95807 239979 95835
rect 240007 95807 240041 95835
rect 240069 95807 256437 95835
rect 256465 95807 256499 95835
rect 256527 95807 256561 95835
rect 256589 95807 256623 95835
rect 256651 95807 265437 95835
rect 265465 95807 265499 95835
rect 265527 95807 265561 95835
rect 265589 95807 265623 95835
rect 265651 95807 274437 95835
rect 274465 95807 274499 95835
rect 274527 95807 274561 95835
rect 274589 95807 274623 95835
rect 274651 95807 283437 95835
rect 283465 95807 283499 95835
rect 283527 95807 283561 95835
rect 283589 95807 283623 95835
rect 283651 95807 292437 95835
rect 292465 95807 292499 95835
rect 292527 95807 292561 95835
rect 292589 95807 292623 95835
rect 292651 95807 299736 95835
rect 299764 95807 299798 95835
rect 299826 95807 299860 95835
rect 299888 95807 299922 95835
rect 299950 95807 299998 95835
rect -6 95773 299998 95807
rect -6 95745 42 95773
rect 70 95745 104 95773
rect 132 95745 166 95773
rect 194 95745 228 95773
rect 256 95745 4437 95773
rect 4465 95745 4499 95773
rect 4527 95745 4561 95773
rect 4589 95745 4623 95773
rect 4651 95745 13437 95773
rect 13465 95745 13499 95773
rect 13527 95745 13561 95773
rect 13589 95745 13623 95773
rect 13651 95745 22437 95773
rect 22465 95745 22499 95773
rect 22527 95745 22561 95773
rect 22589 95745 22623 95773
rect 22651 95745 24939 95773
rect 24967 95745 25001 95773
rect 25029 95745 31437 95773
rect 31465 95745 31499 95773
rect 31527 95745 31561 95773
rect 31589 95745 31623 95773
rect 31651 95745 40299 95773
rect 40327 95745 40361 95773
rect 40389 95745 55659 95773
rect 55687 95745 55721 95773
rect 55749 95745 71019 95773
rect 71047 95745 71081 95773
rect 71109 95745 86379 95773
rect 86407 95745 86441 95773
rect 86469 95745 101739 95773
rect 101767 95745 101801 95773
rect 101829 95745 117099 95773
rect 117127 95745 117161 95773
rect 117189 95745 132459 95773
rect 132487 95745 132521 95773
rect 132549 95745 147819 95773
rect 147847 95745 147881 95773
rect 147909 95745 163179 95773
rect 163207 95745 163241 95773
rect 163269 95745 178539 95773
rect 178567 95745 178601 95773
rect 178629 95745 193899 95773
rect 193927 95745 193961 95773
rect 193989 95745 209259 95773
rect 209287 95745 209321 95773
rect 209349 95745 224619 95773
rect 224647 95745 224681 95773
rect 224709 95745 239979 95773
rect 240007 95745 240041 95773
rect 240069 95745 256437 95773
rect 256465 95745 256499 95773
rect 256527 95745 256561 95773
rect 256589 95745 256623 95773
rect 256651 95745 265437 95773
rect 265465 95745 265499 95773
rect 265527 95745 265561 95773
rect 265589 95745 265623 95773
rect 265651 95745 274437 95773
rect 274465 95745 274499 95773
rect 274527 95745 274561 95773
rect 274589 95745 274623 95773
rect 274651 95745 283437 95773
rect 283465 95745 283499 95773
rect 283527 95745 283561 95773
rect 283589 95745 283623 95773
rect 283651 95745 292437 95773
rect 292465 95745 292499 95773
rect 292527 95745 292561 95773
rect 292589 95745 292623 95773
rect 292651 95745 299736 95773
rect 299764 95745 299798 95773
rect 299826 95745 299860 95773
rect 299888 95745 299922 95773
rect 299950 95745 299998 95773
rect -6 95697 299998 95745
rect -6 92959 299998 93007
rect -6 92931 522 92959
rect 550 92931 584 92959
rect 612 92931 646 92959
rect 674 92931 708 92959
rect 736 92931 2577 92959
rect 2605 92931 2639 92959
rect 2667 92931 2701 92959
rect 2729 92931 2763 92959
rect 2791 92931 11577 92959
rect 11605 92931 11639 92959
rect 11667 92931 11701 92959
rect 11729 92931 11763 92959
rect 11791 92931 17259 92959
rect 17287 92931 17321 92959
rect 17349 92931 20577 92959
rect 20605 92931 20639 92959
rect 20667 92931 20701 92959
rect 20729 92931 20763 92959
rect 20791 92931 29577 92959
rect 29605 92931 29639 92959
rect 29667 92931 29701 92959
rect 29729 92931 29763 92959
rect 29791 92931 32619 92959
rect 32647 92931 32681 92959
rect 32709 92931 47979 92959
rect 48007 92931 48041 92959
rect 48069 92931 63339 92959
rect 63367 92931 63401 92959
rect 63429 92931 78699 92959
rect 78727 92931 78761 92959
rect 78789 92931 94059 92959
rect 94087 92931 94121 92959
rect 94149 92931 109419 92959
rect 109447 92931 109481 92959
rect 109509 92931 124779 92959
rect 124807 92931 124841 92959
rect 124869 92931 140139 92959
rect 140167 92931 140201 92959
rect 140229 92931 155499 92959
rect 155527 92931 155561 92959
rect 155589 92931 170859 92959
rect 170887 92931 170921 92959
rect 170949 92931 186219 92959
rect 186247 92931 186281 92959
rect 186309 92931 201579 92959
rect 201607 92931 201641 92959
rect 201669 92931 216939 92959
rect 216967 92931 217001 92959
rect 217029 92931 232299 92959
rect 232327 92931 232361 92959
rect 232389 92931 247659 92959
rect 247687 92931 247721 92959
rect 247749 92931 254577 92959
rect 254605 92931 254639 92959
rect 254667 92931 254701 92959
rect 254729 92931 254763 92959
rect 254791 92931 263577 92959
rect 263605 92931 263639 92959
rect 263667 92931 263701 92959
rect 263729 92931 263763 92959
rect 263791 92931 272577 92959
rect 272605 92931 272639 92959
rect 272667 92931 272701 92959
rect 272729 92931 272763 92959
rect 272791 92931 281577 92959
rect 281605 92931 281639 92959
rect 281667 92931 281701 92959
rect 281729 92931 281763 92959
rect 281791 92931 290577 92959
rect 290605 92931 290639 92959
rect 290667 92931 290701 92959
rect 290729 92931 290763 92959
rect 290791 92931 299256 92959
rect 299284 92931 299318 92959
rect 299346 92931 299380 92959
rect 299408 92931 299442 92959
rect 299470 92931 299998 92959
rect -6 92897 299998 92931
rect -6 92869 522 92897
rect 550 92869 584 92897
rect 612 92869 646 92897
rect 674 92869 708 92897
rect 736 92869 2577 92897
rect 2605 92869 2639 92897
rect 2667 92869 2701 92897
rect 2729 92869 2763 92897
rect 2791 92869 11577 92897
rect 11605 92869 11639 92897
rect 11667 92869 11701 92897
rect 11729 92869 11763 92897
rect 11791 92869 17259 92897
rect 17287 92869 17321 92897
rect 17349 92869 20577 92897
rect 20605 92869 20639 92897
rect 20667 92869 20701 92897
rect 20729 92869 20763 92897
rect 20791 92869 29577 92897
rect 29605 92869 29639 92897
rect 29667 92869 29701 92897
rect 29729 92869 29763 92897
rect 29791 92869 32619 92897
rect 32647 92869 32681 92897
rect 32709 92869 47979 92897
rect 48007 92869 48041 92897
rect 48069 92869 63339 92897
rect 63367 92869 63401 92897
rect 63429 92869 78699 92897
rect 78727 92869 78761 92897
rect 78789 92869 94059 92897
rect 94087 92869 94121 92897
rect 94149 92869 109419 92897
rect 109447 92869 109481 92897
rect 109509 92869 124779 92897
rect 124807 92869 124841 92897
rect 124869 92869 140139 92897
rect 140167 92869 140201 92897
rect 140229 92869 155499 92897
rect 155527 92869 155561 92897
rect 155589 92869 170859 92897
rect 170887 92869 170921 92897
rect 170949 92869 186219 92897
rect 186247 92869 186281 92897
rect 186309 92869 201579 92897
rect 201607 92869 201641 92897
rect 201669 92869 216939 92897
rect 216967 92869 217001 92897
rect 217029 92869 232299 92897
rect 232327 92869 232361 92897
rect 232389 92869 247659 92897
rect 247687 92869 247721 92897
rect 247749 92869 254577 92897
rect 254605 92869 254639 92897
rect 254667 92869 254701 92897
rect 254729 92869 254763 92897
rect 254791 92869 263577 92897
rect 263605 92869 263639 92897
rect 263667 92869 263701 92897
rect 263729 92869 263763 92897
rect 263791 92869 272577 92897
rect 272605 92869 272639 92897
rect 272667 92869 272701 92897
rect 272729 92869 272763 92897
rect 272791 92869 281577 92897
rect 281605 92869 281639 92897
rect 281667 92869 281701 92897
rect 281729 92869 281763 92897
rect 281791 92869 290577 92897
rect 290605 92869 290639 92897
rect 290667 92869 290701 92897
rect 290729 92869 290763 92897
rect 290791 92869 299256 92897
rect 299284 92869 299318 92897
rect 299346 92869 299380 92897
rect 299408 92869 299442 92897
rect 299470 92869 299998 92897
rect -6 92835 299998 92869
rect -6 92807 522 92835
rect 550 92807 584 92835
rect 612 92807 646 92835
rect 674 92807 708 92835
rect 736 92807 2577 92835
rect 2605 92807 2639 92835
rect 2667 92807 2701 92835
rect 2729 92807 2763 92835
rect 2791 92807 11577 92835
rect 11605 92807 11639 92835
rect 11667 92807 11701 92835
rect 11729 92807 11763 92835
rect 11791 92807 17259 92835
rect 17287 92807 17321 92835
rect 17349 92807 20577 92835
rect 20605 92807 20639 92835
rect 20667 92807 20701 92835
rect 20729 92807 20763 92835
rect 20791 92807 29577 92835
rect 29605 92807 29639 92835
rect 29667 92807 29701 92835
rect 29729 92807 29763 92835
rect 29791 92807 32619 92835
rect 32647 92807 32681 92835
rect 32709 92807 47979 92835
rect 48007 92807 48041 92835
rect 48069 92807 63339 92835
rect 63367 92807 63401 92835
rect 63429 92807 78699 92835
rect 78727 92807 78761 92835
rect 78789 92807 94059 92835
rect 94087 92807 94121 92835
rect 94149 92807 109419 92835
rect 109447 92807 109481 92835
rect 109509 92807 124779 92835
rect 124807 92807 124841 92835
rect 124869 92807 140139 92835
rect 140167 92807 140201 92835
rect 140229 92807 155499 92835
rect 155527 92807 155561 92835
rect 155589 92807 170859 92835
rect 170887 92807 170921 92835
rect 170949 92807 186219 92835
rect 186247 92807 186281 92835
rect 186309 92807 201579 92835
rect 201607 92807 201641 92835
rect 201669 92807 216939 92835
rect 216967 92807 217001 92835
rect 217029 92807 232299 92835
rect 232327 92807 232361 92835
rect 232389 92807 247659 92835
rect 247687 92807 247721 92835
rect 247749 92807 254577 92835
rect 254605 92807 254639 92835
rect 254667 92807 254701 92835
rect 254729 92807 254763 92835
rect 254791 92807 263577 92835
rect 263605 92807 263639 92835
rect 263667 92807 263701 92835
rect 263729 92807 263763 92835
rect 263791 92807 272577 92835
rect 272605 92807 272639 92835
rect 272667 92807 272701 92835
rect 272729 92807 272763 92835
rect 272791 92807 281577 92835
rect 281605 92807 281639 92835
rect 281667 92807 281701 92835
rect 281729 92807 281763 92835
rect 281791 92807 290577 92835
rect 290605 92807 290639 92835
rect 290667 92807 290701 92835
rect 290729 92807 290763 92835
rect 290791 92807 299256 92835
rect 299284 92807 299318 92835
rect 299346 92807 299380 92835
rect 299408 92807 299442 92835
rect 299470 92807 299998 92835
rect -6 92773 299998 92807
rect -6 92745 522 92773
rect 550 92745 584 92773
rect 612 92745 646 92773
rect 674 92745 708 92773
rect 736 92745 2577 92773
rect 2605 92745 2639 92773
rect 2667 92745 2701 92773
rect 2729 92745 2763 92773
rect 2791 92745 11577 92773
rect 11605 92745 11639 92773
rect 11667 92745 11701 92773
rect 11729 92745 11763 92773
rect 11791 92745 17259 92773
rect 17287 92745 17321 92773
rect 17349 92745 20577 92773
rect 20605 92745 20639 92773
rect 20667 92745 20701 92773
rect 20729 92745 20763 92773
rect 20791 92745 29577 92773
rect 29605 92745 29639 92773
rect 29667 92745 29701 92773
rect 29729 92745 29763 92773
rect 29791 92745 32619 92773
rect 32647 92745 32681 92773
rect 32709 92745 47979 92773
rect 48007 92745 48041 92773
rect 48069 92745 63339 92773
rect 63367 92745 63401 92773
rect 63429 92745 78699 92773
rect 78727 92745 78761 92773
rect 78789 92745 94059 92773
rect 94087 92745 94121 92773
rect 94149 92745 109419 92773
rect 109447 92745 109481 92773
rect 109509 92745 124779 92773
rect 124807 92745 124841 92773
rect 124869 92745 140139 92773
rect 140167 92745 140201 92773
rect 140229 92745 155499 92773
rect 155527 92745 155561 92773
rect 155589 92745 170859 92773
rect 170887 92745 170921 92773
rect 170949 92745 186219 92773
rect 186247 92745 186281 92773
rect 186309 92745 201579 92773
rect 201607 92745 201641 92773
rect 201669 92745 216939 92773
rect 216967 92745 217001 92773
rect 217029 92745 232299 92773
rect 232327 92745 232361 92773
rect 232389 92745 247659 92773
rect 247687 92745 247721 92773
rect 247749 92745 254577 92773
rect 254605 92745 254639 92773
rect 254667 92745 254701 92773
rect 254729 92745 254763 92773
rect 254791 92745 263577 92773
rect 263605 92745 263639 92773
rect 263667 92745 263701 92773
rect 263729 92745 263763 92773
rect 263791 92745 272577 92773
rect 272605 92745 272639 92773
rect 272667 92745 272701 92773
rect 272729 92745 272763 92773
rect 272791 92745 281577 92773
rect 281605 92745 281639 92773
rect 281667 92745 281701 92773
rect 281729 92745 281763 92773
rect 281791 92745 290577 92773
rect 290605 92745 290639 92773
rect 290667 92745 290701 92773
rect 290729 92745 290763 92773
rect 290791 92745 299256 92773
rect 299284 92745 299318 92773
rect 299346 92745 299380 92773
rect 299408 92745 299442 92773
rect 299470 92745 299998 92773
rect -6 92697 299998 92745
rect -6 86959 299998 87007
rect -6 86931 42 86959
rect 70 86931 104 86959
rect 132 86931 166 86959
rect 194 86931 228 86959
rect 256 86931 4437 86959
rect 4465 86931 4499 86959
rect 4527 86931 4561 86959
rect 4589 86931 4623 86959
rect 4651 86931 13437 86959
rect 13465 86931 13499 86959
rect 13527 86931 13561 86959
rect 13589 86931 13623 86959
rect 13651 86931 22437 86959
rect 22465 86931 22499 86959
rect 22527 86931 22561 86959
rect 22589 86931 22623 86959
rect 22651 86931 24939 86959
rect 24967 86931 25001 86959
rect 25029 86931 31437 86959
rect 31465 86931 31499 86959
rect 31527 86931 31561 86959
rect 31589 86931 31623 86959
rect 31651 86931 40299 86959
rect 40327 86931 40361 86959
rect 40389 86931 55659 86959
rect 55687 86931 55721 86959
rect 55749 86931 71019 86959
rect 71047 86931 71081 86959
rect 71109 86931 86379 86959
rect 86407 86931 86441 86959
rect 86469 86931 101739 86959
rect 101767 86931 101801 86959
rect 101829 86931 117099 86959
rect 117127 86931 117161 86959
rect 117189 86931 132459 86959
rect 132487 86931 132521 86959
rect 132549 86931 147819 86959
rect 147847 86931 147881 86959
rect 147909 86931 163179 86959
rect 163207 86931 163241 86959
rect 163269 86931 178539 86959
rect 178567 86931 178601 86959
rect 178629 86931 193899 86959
rect 193927 86931 193961 86959
rect 193989 86931 209259 86959
rect 209287 86931 209321 86959
rect 209349 86931 224619 86959
rect 224647 86931 224681 86959
rect 224709 86931 239979 86959
rect 240007 86931 240041 86959
rect 240069 86931 256437 86959
rect 256465 86931 256499 86959
rect 256527 86931 256561 86959
rect 256589 86931 256623 86959
rect 256651 86931 265437 86959
rect 265465 86931 265499 86959
rect 265527 86931 265561 86959
rect 265589 86931 265623 86959
rect 265651 86931 274437 86959
rect 274465 86931 274499 86959
rect 274527 86931 274561 86959
rect 274589 86931 274623 86959
rect 274651 86931 283437 86959
rect 283465 86931 283499 86959
rect 283527 86931 283561 86959
rect 283589 86931 283623 86959
rect 283651 86931 292437 86959
rect 292465 86931 292499 86959
rect 292527 86931 292561 86959
rect 292589 86931 292623 86959
rect 292651 86931 299736 86959
rect 299764 86931 299798 86959
rect 299826 86931 299860 86959
rect 299888 86931 299922 86959
rect 299950 86931 299998 86959
rect -6 86897 299998 86931
rect -6 86869 42 86897
rect 70 86869 104 86897
rect 132 86869 166 86897
rect 194 86869 228 86897
rect 256 86869 4437 86897
rect 4465 86869 4499 86897
rect 4527 86869 4561 86897
rect 4589 86869 4623 86897
rect 4651 86869 13437 86897
rect 13465 86869 13499 86897
rect 13527 86869 13561 86897
rect 13589 86869 13623 86897
rect 13651 86869 22437 86897
rect 22465 86869 22499 86897
rect 22527 86869 22561 86897
rect 22589 86869 22623 86897
rect 22651 86869 24939 86897
rect 24967 86869 25001 86897
rect 25029 86869 31437 86897
rect 31465 86869 31499 86897
rect 31527 86869 31561 86897
rect 31589 86869 31623 86897
rect 31651 86869 40299 86897
rect 40327 86869 40361 86897
rect 40389 86869 55659 86897
rect 55687 86869 55721 86897
rect 55749 86869 71019 86897
rect 71047 86869 71081 86897
rect 71109 86869 86379 86897
rect 86407 86869 86441 86897
rect 86469 86869 101739 86897
rect 101767 86869 101801 86897
rect 101829 86869 117099 86897
rect 117127 86869 117161 86897
rect 117189 86869 132459 86897
rect 132487 86869 132521 86897
rect 132549 86869 147819 86897
rect 147847 86869 147881 86897
rect 147909 86869 163179 86897
rect 163207 86869 163241 86897
rect 163269 86869 178539 86897
rect 178567 86869 178601 86897
rect 178629 86869 193899 86897
rect 193927 86869 193961 86897
rect 193989 86869 209259 86897
rect 209287 86869 209321 86897
rect 209349 86869 224619 86897
rect 224647 86869 224681 86897
rect 224709 86869 239979 86897
rect 240007 86869 240041 86897
rect 240069 86869 256437 86897
rect 256465 86869 256499 86897
rect 256527 86869 256561 86897
rect 256589 86869 256623 86897
rect 256651 86869 265437 86897
rect 265465 86869 265499 86897
rect 265527 86869 265561 86897
rect 265589 86869 265623 86897
rect 265651 86869 274437 86897
rect 274465 86869 274499 86897
rect 274527 86869 274561 86897
rect 274589 86869 274623 86897
rect 274651 86869 283437 86897
rect 283465 86869 283499 86897
rect 283527 86869 283561 86897
rect 283589 86869 283623 86897
rect 283651 86869 292437 86897
rect 292465 86869 292499 86897
rect 292527 86869 292561 86897
rect 292589 86869 292623 86897
rect 292651 86869 299736 86897
rect 299764 86869 299798 86897
rect 299826 86869 299860 86897
rect 299888 86869 299922 86897
rect 299950 86869 299998 86897
rect -6 86835 299998 86869
rect -6 86807 42 86835
rect 70 86807 104 86835
rect 132 86807 166 86835
rect 194 86807 228 86835
rect 256 86807 4437 86835
rect 4465 86807 4499 86835
rect 4527 86807 4561 86835
rect 4589 86807 4623 86835
rect 4651 86807 13437 86835
rect 13465 86807 13499 86835
rect 13527 86807 13561 86835
rect 13589 86807 13623 86835
rect 13651 86807 22437 86835
rect 22465 86807 22499 86835
rect 22527 86807 22561 86835
rect 22589 86807 22623 86835
rect 22651 86807 24939 86835
rect 24967 86807 25001 86835
rect 25029 86807 31437 86835
rect 31465 86807 31499 86835
rect 31527 86807 31561 86835
rect 31589 86807 31623 86835
rect 31651 86807 40299 86835
rect 40327 86807 40361 86835
rect 40389 86807 55659 86835
rect 55687 86807 55721 86835
rect 55749 86807 71019 86835
rect 71047 86807 71081 86835
rect 71109 86807 86379 86835
rect 86407 86807 86441 86835
rect 86469 86807 101739 86835
rect 101767 86807 101801 86835
rect 101829 86807 117099 86835
rect 117127 86807 117161 86835
rect 117189 86807 132459 86835
rect 132487 86807 132521 86835
rect 132549 86807 147819 86835
rect 147847 86807 147881 86835
rect 147909 86807 163179 86835
rect 163207 86807 163241 86835
rect 163269 86807 178539 86835
rect 178567 86807 178601 86835
rect 178629 86807 193899 86835
rect 193927 86807 193961 86835
rect 193989 86807 209259 86835
rect 209287 86807 209321 86835
rect 209349 86807 224619 86835
rect 224647 86807 224681 86835
rect 224709 86807 239979 86835
rect 240007 86807 240041 86835
rect 240069 86807 256437 86835
rect 256465 86807 256499 86835
rect 256527 86807 256561 86835
rect 256589 86807 256623 86835
rect 256651 86807 265437 86835
rect 265465 86807 265499 86835
rect 265527 86807 265561 86835
rect 265589 86807 265623 86835
rect 265651 86807 274437 86835
rect 274465 86807 274499 86835
rect 274527 86807 274561 86835
rect 274589 86807 274623 86835
rect 274651 86807 283437 86835
rect 283465 86807 283499 86835
rect 283527 86807 283561 86835
rect 283589 86807 283623 86835
rect 283651 86807 292437 86835
rect 292465 86807 292499 86835
rect 292527 86807 292561 86835
rect 292589 86807 292623 86835
rect 292651 86807 299736 86835
rect 299764 86807 299798 86835
rect 299826 86807 299860 86835
rect 299888 86807 299922 86835
rect 299950 86807 299998 86835
rect -6 86773 299998 86807
rect -6 86745 42 86773
rect 70 86745 104 86773
rect 132 86745 166 86773
rect 194 86745 228 86773
rect 256 86745 4437 86773
rect 4465 86745 4499 86773
rect 4527 86745 4561 86773
rect 4589 86745 4623 86773
rect 4651 86745 13437 86773
rect 13465 86745 13499 86773
rect 13527 86745 13561 86773
rect 13589 86745 13623 86773
rect 13651 86745 22437 86773
rect 22465 86745 22499 86773
rect 22527 86745 22561 86773
rect 22589 86745 22623 86773
rect 22651 86745 24939 86773
rect 24967 86745 25001 86773
rect 25029 86745 31437 86773
rect 31465 86745 31499 86773
rect 31527 86745 31561 86773
rect 31589 86745 31623 86773
rect 31651 86745 40299 86773
rect 40327 86745 40361 86773
rect 40389 86745 55659 86773
rect 55687 86745 55721 86773
rect 55749 86745 71019 86773
rect 71047 86745 71081 86773
rect 71109 86745 86379 86773
rect 86407 86745 86441 86773
rect 86469 86745 101739 86773
rect 101767 86745 101801 86773
rect 101829 86745 117099 86773
rect 117127 86745 117161 86773
rect 117189 86745 132459 86773
rect 132487 86745 132521 86773
rect 132549 86745 147819 86773
rect 147847 86745 147881 86773
rect 147909 86745 163179 86773
rect 163207 86745 163241 86773
rect 163269 86745 178539 86773
rect 178567 86745 178601 86773
rect 178629 86745 193899 86773
rect 193927 86745 193961 86773
rect 193989 86745 209259 86773
rect 209287 86745 209321 86773
rect 209349 86745 224619 86773
rect 224647 86745 224681 86773
rect 224709 86745 239979 86773
rect 240007 86745 240041 86773
rect 240069 86745 256437 86773
rect 256465 86745 256499 86773
rect 256527 86745 256561 86773
rect 256589 86745 256623 86773
rect 256651 86745 265437 86773
rect 265465 86745 265499 86773
rect 265527 86745 265561 86773
rect 265589 86745 265623 86773
rect 265651 86745 274437 86773
rect 274465 86745 274499 86773
rect 274527 86745 274561 86773
rect 274589 86745 274623 86773
rect 274651 86745 283437 86773
rect 283465 86745 283499 86773
rect 283527 86745 283561 86773
rect 283589 86745 283623 86773
rect 283651 86745 292437 86773
rect 292465 86745 292499 86773
rect 292527 86745 292561 86773
rect 292589 86745 292623 86773
rect 292651 86745 299736 86773
rect 299764 86745 299798 86773
rect 299826 86745 299860 86773
rect 299888 86745 299922 86773
rect 299950 86745 299998 86773
rect -6 86697 299998 86745
rect -6 83959 299998 84007
rect -6 83931 522 83959
rect 550 83931 584 83959
rect 612 83931 646 83959
rect 674 83931 708 83959
rect 736 83931 2577 83959
rect 2605 83931 2639 83959
rect 2667 83931 2701 83959
rect 2729 83931 2763 83959
rect 2791 83931 11577 83959
rect 11605 83931 11639 83959
rect 11667 83931 11701 83959
rect 11729 83931 11763 83959
rect 11791 83931 17259 83959
rect 17287 83931 17321 83959
rect 17349 83931 20577 83959
rect 20605 83931 20639 83959
rect 20667 83931 20701 83959
rect 20729 83931 20763 83959
rect 20791 83931 29577 83959
rect 29605 83931 29639 83959
rect 29667 83931 29701 83959
rect 29729 83931 29763 83959
rect 29791 83931 32619 83959
rect 32647 83931 32681 83959
rect 32709 83931 47979 83959
rect 48007 83931 48041 83959
rect 48069 83931 63339 83959
rect 63367 83931 63401 83959
rect 63429 83931 78699 83959
rect 78727 83931 78761 83959
rect 78789 83931 94059 83959
rect 94087 83931 94121 83959
rect 94149 83931 109419 83959
rect 109447 83931 109481 83959
rect 109509 83931 124779 83959
rect 124807 83931 124841 83959
rect 124869 83931 140139 83959
rect 140167 83931 140201 83959
rect 140229 83931 155499 83959
rect 155527 83931 155561 83959
rect 155589 83931 170859 83959
rect 170887 83931 170921 83959
rect 170949 83931 186219 83959
rect 186247 83931 186281 83959
rect 186309 83931 201579 83959
rect 201607 83931 201641 83959
rect 201669 83931 216939 83959
rect 216967 83931 217001 83959
rect 217029 83931 232299 83959
rect 232327 83931 232361 83959
rect 232389 83931 247659 83959
rect 247687 83931 247721 83959
rect 247749 83931 254577 83959
rect 254605 83931 254639 83959
rect 254667 83931 254701 83959
rect 254729 83931 254763 83959
rect 254791 83931 263577 83959
rect 263605 83931 263639 83959
rect 263667 83931 263701 83959
rect 263729 83931 263763 83959
rect 263791 83931 272577 83959
rect 272605 83931 272639 83959
rect 272667 83931 272701 83959
rect 272729 83931 272763 83959
rect 272791 83931 281577 83959
rect 281605 83931 281639 83959
rect 281667 83931 281701 83959
rect 281729 83931 281763 83959
rect 281791 83931 290577 83959
rect 290605 83931 290639 83959
rect 290667 83931 290701 83959
rect 290729 83931 290763 83959
rect 290791 83931 299256 83959
rect 299284 83931 299318 83959
rect 299346 83931 299380 83959
rect 299408 83931 299442 83959
rect 299470 83931 299998 83959
rect -6 83897 299998 83931
rect -6 83869 522 83897
rect 550 83869 584 83897
rect 612 83869 646 83897
rect 674 83869 708 83897
rect 736 83869 2577 83897
rect 2605 83869 2639 83897
rect 2667 83869 2701 83897
rect 2729 83869 2763 83897
rect 2791 83869 11577 83897
rect 11605 83869 11639 83897
rect 11667 83869 11701 83897
rect 11729 83869 11763 83897
rect 11791 83869 17259 83897
rect 17287 83869 17321 83897
rect 17349 83869 20577 83897
rect 20605 83869 20639 83897
rect 20667 83869 20701 83897
rect 20729 83869 20763 83897
rect 20791 83869 29577 83897
rect 29605 83869 29639 83897
rect 29667 83869 29701 83897
rect 29729 83869 29763 83897
rect 29791 83869 32619 83897
rect 32647 83869 32681 83897
rect 32709 83869 47979 83897
rect 48007 83869 48041 83897
rect 48069 83869 63339 83897
rect 63367 83869 63401 83897
rect 63429 83869 78699 83897
rect 78727 83869 78761 83897
rect 78789 83869 94059 83897
rect 94087 83869 94121 83897
rect 94149 83869 109419 83897
rect 109447 83869 109481 83897
rect 109509 83869 124779 83897
rect 124807 83869 124841 83897
rect 124869 83869 140139 83897
rect 140167 83869 140201 83897
rect 140229 83869 155499 83897
rect 155527 83869 155561 83897
rect 155589 83869 170859 83897
rect 170887 83869 170921 83897
rect 170949 83869 186219 83897
rect 186247 83869 186281 83897
rect 186309 83869 201579 83897
rect 201607 83869 201641 83897
rect 201669 83869 216939 83897
rect 216967 83869 217001 83897
rect 217029 83869 232299 83897
rect 232327 83869 232361 83897
rect 232389 83869 247659 83897
rect 247687 83869 247721 83897
rect 247749 83869 254577 83897
rect 254605 83869 254639 83897
rect 254667 83869 254701 83897
rect 254729 83869 254763 83897
rect 254791 83869 263577 83897
rect 263605 83869 263639 83897
rect 263667 83869 263701 83897
rect 263729 83869 263763 83897
rect 263791 83869 272577 83897
rect 272605 83869 272639 83897
rect 272667 83869 272701 83897
rect 272729 83869 272763 83897
rect 272791 83869 281577 83897
rect 281605 83869 281639 83897
rect 281667 83869 281701 83897
rect 281729 83869 281763 83897
rect 281791 83869 290577 83897
rect 290605 83869 290639 83897
rect 290667 83869 290701 83897
rect 290729 83869 290763 83897
rect 290791 83869 299256 83897
rect 299284 83869 299318 83897
rect 299346 83869 299380 83897
rect 299408 83869 299442 83897
rect 299470 83869 299998 83897
rect -6 83835 299998 83869
rect -6 83807 522 83835
rect 550 83807 584 83835
rect 612 83807 646 83835
rect 674 83807 708 83835
rect 736 83807 2577 83835
rect 2605 83807 2639 83835
rect 2667 83807 2701 83835
rect 2729 83807 2763 83835
rect 2791 83807 11577 83835
rect 11605 83807 11639 83835
rect 11667 83807 11701 83835
rect 11729 83807 11763 83835
rect 11791 83807 17259 83835
rect 17287 83807 17321 83835
rect 17349 83807 20577 83835
rect 20605 83807 20639 83835
rect 20667 83807 20701 83835
rect 20729 83807 20763 83835
rect 20791 83807 29577 83835
rect 29605 83807 29639 83835
rect 29667 83807 29701 83835
rect 29729 83807 29763 83835
rect 29791 83807 32619 83835
rect 32647 83807 32681 83835
rect 32709 83807 47979 83835
rect 48007 83807 48041 83835
rect 48069 83807 63339 83835
rect 63367 83807 63401 83835
rect 63429 83807 78699 83835
rect 78727 83807 78761 83835
rect 78789 83807 94059 83835
rect 94087 83807 94121 83835
rect 94149 83807 109419 83835
rect 109447 83807 109481 83835
rect 109509 83807 124779 83835
rect 124807 83807 124841 83835
rect 124869 83807 140139 83835
rect 140167 83807 140201 83835
rect 140229 83807 155499 83835
rect 155527 83807 155561 83835
rect 155589 83807 170859 83835
rect 170887 83807 170921 83835
rect 170949 83807 186219 83835
rect 186247 83807 186281 83835
rect 186309 83807 201579 83835
rect 201607 83807 201641 83835
rect 201669 83807 216939 83835
rect 216967 83807 217001 83835
rect 217029 83807 232299 83835
rect 232327 83807 232361 83835
rect 232389 83807 247659 83835
rect 247687 83807 247721 83835
rect 247749 83807 254577 83835
rect 254605 83807 254639 83835
rect 254667 83807 254701 83835
rect 254729 83807 254763 83835
rect 254791 83807 263577 83835
rect 263605 83807 263639 83835
rect 263667 83807 263701 83835
rect 263729 83807 263763 83835
rect 263791 83807 272577 83835
rect 272605 83807 272639 83835
rect 272667 83807 272701 83835
rect 272729 83807 272763 83835
rect 272791 83807 281577 83835
rect 281605 83807 281639 83835
rect 281667 83807 281701 83835
rect 281729 83807 281763 83835
rect 281791 83807 290577 83835
rect 290605 83807 290639 83835
rect 290667 83807 290701 83835
rect 290729 83807 290763 83835
rect 290791 83807 299256 83835
rect 299284 83807 299318 83835
rect 299346 83807 299380 83835
rect 299408 83807 299442 83835
rect 299470 83807 299998 83835
rect -6 83773 299998 83807
rect -6 83745 522 83773
rect 550 83745 584 83773
rect 612 83745 646 83773
rect 674 83745 708 83773
rect 736 83745 2577 83773
rect 2605 83745 2639 83773
rect 2667 83745 2701 83773
rect 2729 83745 2763 83773
rect 2791 83745 11577 83773
rect 11605 83745 11639 83773
rect 11667 83745 11701 83773
rect 11729 83745 11763 83773
rect 11791 83745 17259 83773
rect 17287 83745 17321 83773
rect 17349 83745 20577 83773
rect 20605 83745 20639 83773
rect 20667 83745 20701 83773
rect 20729 83745 20763 83773
rect 20791 83745 29577 83773
rect 29605 83745 29639 83773
rect 29667 83745 29701 83773
rect 29729 83745 29763 83773
rect 29791 83745 32619 83773
rect 32647 83745 32681 83773
rect 32709 83745 47979 83773
rect 48007 83745 48041 83773
rect 48069 83745 63339 83773
rect 63367 83745 63401 83773
rect 63429 83745 78699 83773
rect 78727 83745 78761 83773
rect 78789 83745 94059 83773
rect 94087 83745 94121 83773
rect 94149 83745 109419 83773
rect 109447 83745 109481 83773
rect 109509 83745 124779 83773
rect 124807 83745 124841 83773
rect 124869 83745 140139 83773
rect 140167 83745 140201 83773
rect 140229 83745 155499 83773
rect 155527 83745 155561 83773
rect 155589 83745 170859 83773
rect 170887 83745 170921 83773
rect 170949 83745 186219 83773
rect 186247 83745 186281 83773
rect 186309 83745 201579 83773
rect 201607 83745 201641 83773
rect 201669 83745 216939 83773
rect 216967 83745 217001 83773
rect 217029 83745 232299 83773
rect 232327 83745 232361 83773
rect 232389 83745 247659 83773
rect 247687 83745 247721 83773
rect 247749 83745 254577 83773
rect 254605 83745 254639 83773
rect 254667 83745 254701 83773
rect 254729 83745 254763 83773
rect 254791 83745 263577 83773
rect 263605 83745 263639 83773
rect 263667 83745 263701 83773
rect 263729 83745 263763 83773
rect 263791 83745 272577 83773
rect 272605 83745 272639 83773
rect 272667 83745 272701 83773
rect 272729 83745 272763 83773
rect 272791 83745 281577 83773
rect 281605 83745 281639 83773
rect 281667 83745 281701 83773
rect 281729 83745 281763 83773
rect 281791 83745 290577 83773
rect 290605 83745 290639 83773
rect 290667 83745 290701 83773
rect 290729 83745 290763 83773
rect 290791 83745 299256 83773
rect 299284 83745 299318 83773
rect 299346 83745 299380 83773
rect 299408 83745 299442 83773
rect 299470 83745 299998 83773
rect -6 83697 299998 83745
rect -6 77959 299998 78007
rect -6 77931 42 77959
rect 70 77931 104 77959
rect 132 77931 166 77959
rect 194 77931 228 77959
rect 256 77931 4437 77959
rect 4465 77931 4499 77959
rect 4527 77931 4561 77959
rect 4589 77931 4623 77959
rect 4651 77931 13437 77959
rect 13465 77931 13499 77959
rect 13527 77931 13561 77959
rect 13589 77931 13623 77959
rect 13651 77931 22437 77959
rect 22465 77931 22499 77959
rect 22527 77931 22561 77959
rect 22589 77931 22623 77959
rect 22651 77931 24939 77959
rect 24967 77931 25001 77959
rect 25029 77931 31437 77959
rect 31465 77931 31499 77959
rect 31527 77931 31561 77959
rect 31589 77931 31623 77959
rect 31651 77931 40299 77959
rect 40327 77931 40361 77959
rect 40389 77931 55659 77959
rect 55687 77931 55721 77959
rect 55749 77931 71019 77959
rect 71047 77931 71081 77959
rect 71109 77931 86379 77959
rect 86407 77931 86441 77959
rect 86469 77931 101739 77959
rect 101767 77931 101801 77959
rect 101829 77931 117099 77959
rect 117127 77931 117161 77959
rect 117189 77931 132459 77959
rect 132487 77931 132521 77959
rect 132549 77931 147819 77959
rect 147847 77931 147881 77959
rect 147909 77931 163179 77959
rect 163207 77931 163241 77959
rect 163269 77931 178539 77959
rect 178567 77931 178601 77959
rect 178629 77931 193899 77959
rect 193927 77931 193961 77959
rect 193989 77931 209259 77959
rect 209287 77931 209321 77959
rect 209349 77931 224619 77959
rect 224647 77931 224681 77959
rect 224709 77931 239979 77959
rect 240007 77931 240041 77959
rect 240069 77931 256437 77959
rect 256465 77931 256499 77959
rect 256527 77931 256561 77959
rect 256589 77931 256623 77959
rect 256651 77931 265437 77959
rect 265465 77931 265499 77959
rect 265527 77931 265561 77959
rect 265589 77931 265623 77959
rect 265651 77931 274437 77959
rect 274465 77931 274499 77959
rect 274527 77931 274561 77959
rect 274589 77931 274623 77959
rect 274651 77931 283437 77959
rect 283465 77931 283499 77959
rect 283527 77931 283561 77959
rect 283589 77931 283623 77959
rect 283651 77931 292437 77959
rect 292465 77931 292499 77959
rect 292527 77931 292561 77959
rect 292589 77931 292623 77959
rect 292651 77931 299736 77959
rect 299764 77931 299798 77959
rect 299826 77931 299860 77959
rect 299888 77931 299922 77959
rect 299950 77931 299998 77959
rect -6 77897 299998 77931
rect -6 77869 42 77897
rect 70 77869 104 77897
rect 132 77869 166 77897
rect 194 77869 228 77897
rect 256 77869 4437 77897
rect 4465 77869 4499 77897
rect 4527 77869 4561 77897
rect 4589 77869 4623 77897
rect 4651 77869 13437 77897
rect 13465 77869 13499 77897
rect 13527 77869 13561 77897
rect 13589 77869 13623 77897
rect 13651 77869 22437 77897
rect 22465 77869 22499 77897
rect 22527 77869 22561 77897
rect 22589 77869 22623 77897
rect 22651 77869 24939 77897
rect 24967 77869 25001 77897
rect 25029 77869 31437 77897
rect 31465 77869 31499 77897
rect 31527 77869 31561 77897
rect 31589 77869 31623 77897
rect 31651 77869 40299 77897
rect 40327 77869 40361 77897
rect 40389 77869 55659 77897
rect 55687 77869 55721 77897
rect 55749 77869 71019 77897
rect 71047 77869 71081 77897
rect 71109 77869 86379 77897
rect 86407 77869 86441 77897
rect 86469 77869 101739 77897
rect 101767 77869 101801 77897
rect 101829 77869 117099 77897
rect 117127 77869 117161 77897
rect 117189 77869 132459 77897
rect 132487 77869 132521 77897
rect 132549 77869 147819 77897
rect 147847 77869 147881 77897
rect 147909 77869 163179 77897
rect 163207 77869 163241 77897
rect 163269 77869 178539 77897
rect 178567 77869 178601 77897
rect 178629 77869 193899 77897
rect 193927 77869 193961 77897
rect 193989 77869 209259 77897
rect 209287 77869 209321 77897
rect 209349 77869 224619 77897
rect 224647 77869 224681 77897
rect 224709 77869 239979 77897
rect 240007 77869 240041 77897
rect 240069 77869 256437 77897
rect 256465 77869 256499 77897
rect 256527 77869 256561 77897
rect 256589 77869 256623 77897
rect 256651 77869 265437 77897
rect 265465 77869 265499 77897
rect 265527 77869 265561 77897
rect 265589 77869 265623 77897
rect 265651 77869 274437 77897
rect 274465 77869 274499 77897
rect 274527 77869 274561 77897
rect 274589 77869 274623 77897
rect 274651 77869 283437 77897
rect 283465 77869 283499 77897
rect 283527 77869 283561 77897
rect 283589 77869 283623 77897
rect 283651 77869 292437 77897
rect 292465 77869 292499 77897
rect 292527 77869 292561 77897
rect 292589 77869 292623 77897
rect 292651 77869 299736 77897
rect 299764 77869 299798 77897
rect 299826 77869 299860 77897
rect 299888 77869 299922 77897
rect 299950 77869 299998 77897
rect -6 77835 299998 77869
rect -6 77807 42 77835
rect 70 77807 104 77835
rect 132 77807 166 77835
rect 194 77807 228 77835
rect 256 77807 4437 77835
rect 4465 77807 4499 77835
rect 4527 77807 4561 77835
rect 4589 77807 4623 77835
rect 4651 77807 13437 77835
rect 13465 77807 13499 77835
rect 13527 77807 13561 77835
rect 13589 77807 13623 77835
rect 13651 77807 22437 77835
rect 22465 77807 22499 77835
rect 22527 77807 22561 77835
rect 22589 77807 22623 77835
rect 22651 77807 24939 77835
rect 24967 77807 25001 77835
rect 25029 77807 31437 77835
rect 31465 77807 31499 77835
rect 31527 77807 31561 77835
rect 31589 77807 31623 77835
rect 31651 77807 40299 77835
rect 40327 77807 40361 77835
rect 40389 77807 55659 77835
rect 55687 77807 55721 77835
rect 55749 77807 71019 77835
rect 71047 77807 71081 77835
rect 71109 77807 86379 77835
rect 86407 77807 86441 77835
rect 86469 77807 101739 77835
rect 101767 77807 101801 77835
rect 101829 77807 117099 77835
rect 117127 77807 117161 77835
rect 117189 77807 132459 77835
rect 132487 77807 132521 77835
rect 132549 77807 147819 77835
rect 147847 77807 147881 77835
rect 147909 77807 163179 77835
rect 163207 77807 163241 77835
rect 163269 77807 178539 77835
rect 178567 77807 178601 77835
rect 178629 77807 193899 77835
rect 193927 77807 193961 77835
rect 193989 77807 209259 77835
rect 209287 77807 209321 77835
rect 209349 77807 224619 77835
rect 224647 77807 224681 77835
rect 224709 77807 239979 77835
rect 240007 77807 240041 77835
rect 240069 77807 256437 77835
rect 256465 77807 256499 77835
rect 256527 77807 256561 77835
rect 256589 77807 256623 77835
rect 256651 77807 265437 77835
rect 265465 77807 265499 77835
rect 265527 77807 265561 77835
rect 265589 77807 265623 77835
rect 265651 77807 274437 77835
rect 274465 77807 274499 77835
rect 274527 77807 274561 77835
rect 274589 77807 274623 77835
rect 274651 77807 283437 77835
rect 283465 77807 283499 77835
rect 283527 77807 283561 77835
rect 283589 77807 283623 77835
rect 283651 77807 292437 77835
rect 292465 77807 292499 77835
rect 292527 77807 292561 77835
rect 292589 77807 292623 77835
rect 292651 77807 299736 77835
rect 299764 77807 299798 77835
rect 299826 77807 299860 77835
rect 299888 77807 299922 77835
rect 299950 77807 299998 77835
rect -6 77773 299998 77807
rect -6 77745 42 77773
rect 70 77745 104 77773
rect 132 77745 166 77773
rect 194 77745 228 77773
rect 256 77745 4437 77773
rect 4465 77745 4499 77773
rect 4527 77745 4561 77773
rect 4589 77745 4623 77773
rect 4651 77745 13437 77773
rect 13465 77745 13499 77773
rect 13527 77745 13561 77773
rect 13589 77745 13623 77773
rect 13651 77745 22437 77773
rect 22465 77745 22499 77773
rect 22527 77745 22561 77773
rect 22589 77745 22623 77773
rect 22651 77745 24939 77773
rect 24967 77745 25001 77773
rect 25029 77745 31437 77773
rect 31465 77745 31499 77773
rect 31527 77745 31561 77773
rect 31589 77745 31623 77773
rect 31651 77745 40299 77773
rect 40327 77745 40361 77773
rect 40389 77745 55659 77773
rect 55687 77745 55721 77773
rect 55749 77745 71019 77773
rect 71047 77745 71081 77773
rect 71109 77745 86379 77773
rect 86407 77745 86441 77773
rect 86469 77745 101739 77773
rect 101767 77745 101801 77773
rect 101829 77745 117099 77773
rect 117127 77745 117161 77773
rect 117189 77745 132459 77773
rect 132487 77745 132521 77773
rect 132549 77745 147819 77773
rect 147847 77745 147881 77773
rect 147909 77745 163179 77773
rect 163207 77745 163241 77773
rect 163269 77745 178539 77773
rect 178567 77745 178601 77773
rect 178629 77745 193899 77773
rect 193927 77745 193961 77773
rect 193989 77745 209259 77773
rect 209287 77745 209321 77773
rect 209349 77745 224619 77773
rect 224647 77745 224681 77773
rect 224709 77745 239979 77773
rect 240007 77745 240041 77773
rect 240069 77745 256437 77773
rect 256465 77745 256499 77773
rect 256527 77745 256561 77773
rect 256589 77745 256623 77773
rect 256651 77745 265437 77773
rect 265465 77745 265499 77773
rect 265527 77745 265561 77773
rect 265589 77745 265623 77773
rect 265651 77745 274437 77773
rect 274465 77745 274499 77773
rect 274527 77745 274561 77773
rect 274589 77745 274623 77773
rect 274651 77745 283437 77773
rect 283465 77745 283499 77773
rect 283527 77745 283561 77773
rect 283589 77745 283623 77773
rect 283651 77745 292437 77773
rect 292465 77745 292499 77773
rect 292527 77745 292561 77773
rect 292589 77745 292623 77773
rect 292651 77745 299736 77773
rect 299764 77745 299798 77773
rect 299826 77745 299860 77773
rect 299888 77745 299922 77773
rect 299950 77745 299998 77773
rect -6 77697 299998 77745
rect -6 74959 299998 75007
rect -6 74931 522 74959
rect 550 74931 584 74959
rect 612 74931 646 74959
rect 674 74931 708 74959
rect 736 74931 2577 74959
rect 2605 74931 2639 74959
rect 2667 74931 2701 74959
rect 2729 74931 2763 74959
rect 2791 74931 11577 74959
rect 11605 74931 11639 74959
rect 11667 74931 11701 74959
rect 11729 74931 11763 74959
rect 11791 74931 17259 74959
rect 17287 74931 17321 74959
rect 17349 74931 20577 74959
rect 20605 74931 20639 74959
rect 20667 74931 20701 74959
rect 20729 74931 20763 74959
rect 20791 74931 29577 74959
rect 29605 74931 29639 74959
rect 29667 74931 29701 74959
rect 29729 74931 29763 74959
rect 29791 74931 32619 74959
rect 32647 74931 32681 74959
rect 32709 74931 47979 74959
rect 48007 74931 48041 74959
rect 48069 74931 63339 74959
rect 63367 74931 63401 74959
rect 63429 74931 78699 74959
rect 78727 74931 78761 74959
rect 78789 74931 94059 74959
rect 94087 74931 94121 74959
rect 94149 74931 109419 74959
rect 109447 74931 109481 74959
rect 109509 74931 124779 74959
rect 124807 74931 124841 74959
rect 124869 74931 140139 74959
rect 140167 74931 140201 74959
rect 140229 74931 155499 74959
rect 155527 74931 155561 74959
rect 155589 74931 170859 74959
rect 170887 74931 170921 74959
rect 170949 74931 186219 74959
rect 186247 74931 186281 74959
rect 186309 74931 201579 74959
rect 201607 74931 201641 74959
rect 201669 74931 216939 74959
rect 216967 74931 217001 74959
rect 217029 74931 232299 74959
rect 232327 74931 232361 74959
rect 232389 74931 247659 74959
rect 247687 74931 247721 74959
rect 247749 74931 254577 74959
rect 254605 74931 254639 74959
rect 254667 74931 254701 74959
rect 254729 74931 254763 74959
rect 254791 74931 263577 74959
rect 263605 74931 263639 74959
rect 263667 74931 263701 74959
rect 263729 74931 263763 74959
rect 263791 74931 272577 74959
rect 272605 74931 272639 74959
rect 272667 74931 272701 74959
rect 272729 74931 272763 74959
rect 272791 74931 281577 74959
rect 281605 74931 281639 74959
rect 281667 74931 281701 74959
rect 281729 74931 281763 74959
rect 281791 74931 290577 74959
rect 290605 74931 290639 74959
rect 290667 74931 290701 74959
rect 290729 74931 290763 74959
rect 290791 74931 299256 74959
rect 299284 74931 299318 74959
rect 299346 74931 299380 74959
rect 299408 74931 299442 74959
rect 299470 74931 299998 74959
rect -6 74897 299998 74931
rect -6 74869 522 74897
rect 550 74869 584 74897
rect 612 74869 646 74897
rect 674 74869 708 74897
rect 736 74869 2577 74897
rect 2605 74869 2639 74897
rect 2667 74869 2701 74897
rect 2729 74869 2763 74897
rect 2791 74869 11577 74897
rect 11605 74869 11639 74897
rect 11667 74869 11701 74897
rect 11729 74869 11763 74897
rect 11791 74869 17259 74897
rect 17287 74869 17321 74897
rect 17349 74869 20577 74897
rect 20605 74869 20639 74897
rect 20667 74869 20701 74897
rect 20729 74869 20763 74897
rect 20791 74869 29577 74897
rect 29605 74869 29639 74897
rect 29667 74869 29701 74897
rect 29729 74869 29763 74897
rect 29791 74869 32619 74897
rect 32647 74869 32681 74897
rect 32709 74869 47979 74897
rect 48007 74869 48041 74897
rect 48069 74869 63339 74897
rect 63367 74869 63401 74897
rect 63429 74869 78699 74897
rect 78727 74869 78761 74897
rect 78789 74869 94059 74897
rect 94087 74869 94121 74897
rect 94149 74869 109419 74897
rect 109447 74869 109481 74897
rect 109509 74869 124779 74897
rect 124807 74869 124841 74897
rect 124869 74869 140139 74897
rect 140167 74869 140201 74897
rect 140229 74869 155499 74897
rect 155527 74869 155561 74897
rect 155589 74869 170859 74897
rect 170887 74869 170921 74897
rect 170949 74869 186219 74897
rect 186247 74869 186281 74897
rect 186309 74869 201579 74897
rect 201607 74869 201641 74897
rect 201669 74869 216939 74897
rect 216967 74869 217001 74897
rect 217029 74869 232299 74897
rect 232327 74869 232361 74897
rect 232389 74869 247659 74897
rect 247687 74869 247721 74897
rect 247749 74869 254577 74897
rect 254605 74869 254639 74897
rect 254667 74869 254701 74897
rect 254729 74869 254763 74897
rect 254791 74869 263577 74897
rect 263605 74869 263639 74897
rect 263667 74869 263701 74897
rect 263729 74869 263763 74897
rect 263791 74869 272577 74897
rect 272605 74869 272639 74897
rect 272667 74869 272701 74897
rect 272729 74869 272763 74897
rect 272791 74869 281577 74897
rect 281605 74869 281639 74897
rect 281667 74869 281701 74897
rect 281729 74869 281763 74897
rect 281791 74869 290577 74897
rect 290605 74869 290639 74897
rect 290667 74869 290701 74897
rect 290729 74869 290763 74897
rect 290791 74869 299256 74897
rect 299284 74869 299318 74897
rect 299346 74869 299380 74897
rect 299408 74869 299442 74897
rect 299470 74869 299998 74897
rect -6 74835 299998 74869
rect -6 74807 522 74835
rect 550 74807 584 74835
rect 612 74807 646 74835
rect 674 74807 708 74835
rect 736 74807 2577 74835
rect 2605 74807 2639 74835
rect 2667 74807 2701 74835
rect 2729 74807 2763 74835
rect 2791 74807 11577 74835
rect 11605 74807 11639 74835
rect 11667 74807 11701 74835
rect 11729 74807 11763 74835
rect 11791 74807 17259 74835
rect 17287 74807 17321 74835
rect 17349 74807 20577 74835
rect 20605 74807 20639 74835
rect 20667 74807 20701 74835
rect 20729 74807 20763 74835
rect 20791 74807 29577 74835
rect 29605 74807 29639 74835
rect 29667 74807 29701 74835
rect 29729 74807 29763 74835
rect 29791 74807 32619 74835
rect 32647 74807 32681 74835
rect 32709 74807 47979 74835
rect 48007 74807 48041 74835
rect 48069 74807 63339 74835
rect 63367 74807 63401 74835
rect 63429 74807 78699 74835
rect 78727 74807 78761 74835
rect 78789 74807 94059 74835
rect 94087 74807 94121 74835
rect 94149 74807 109419 74835
rect 109447 74807 109481 74835
rect 109509 74807 124779 74835
rect 124807 74807 124841 74835
rect 124869 74807 140139 74835
rect 140167 74807 140201 74835
rect 140229 74807 155499 74835
rect 155527 74807 155561 74835
rect 155589 74807 170859 74835
rect 170887 74807 170921 74835
rect 170949 74807 186219 74835
rect 186247 74807 186281 74835
rect 186309 74807 201579 74835
rect 201607 74807 201641 74835
rect 201669 74807 216939 74835
rect 216967 74807 217001 74835
rect 217029 74807 232299 74835
rect 232327 74807 232361 74835
rect 232389 74807 247659 74835
rect 247687 74807 247721 74835
rect 247749 74807 254577 74835
rect 254605 74807 254639 74835
rect 254667 74807 254701 74835
rect 254729 74807 254763 74835
rect 254791 74807 263577 74835
rect 263605 74807 263639 74835
rect 263667 74807 263701 74835
rect 263729 74807 263763 74835
rect 263791 74807 272577 74835
rect 272605 74807 272639 74835
rect 272667 74807 272701 74835
rect 272729 74807 272763 74835
rect 272791 74807 281577 74835
rect 281605 74807 281639 74835
rect 281667 74807 281701 74835
rect 281729 74807 281763 74835
rect 281791 74807 290577 74835
rect 290605 74807 290639 74835
rect 290667 74807 290701 74835
rect 290729 74807 290763 74835
rect 290791 74807 299256 74835
rect 299284 74807 299318 74835
rect 299346 74807 299380 74835
rect 299408 74807 299442 74835
rect 299470 74807 299998 74835
rect -6 74773 299998 74807
rect -6 74745 522 74773
rect 550 74745 584 74773
rect 612 74745 646 74773
rect 674 74745 708 74773
rect 736 74745 2577 74773
rect 2605 74745 2639 74773
rect 2667 74745 2701 74773
rect 2729 74745 2763 74773
rect 2791 74745 11577 74773
rect 11605 74745 11639 74773
rect 11667 74745 11701 74773
rect 11729 74745 11763 74773
rect 11791 74745 17259 74773
rect 17287 74745 17321 74773
rect 17349 74745 20577 74773
rect 20605 74745 20639 74773
rect 20667 74745 20701 74773
rect 20729 74745 20763 74773
rect 20791 74745 29577 74773
rect 29605 74745 29639 74773
rect 29667 74745 29701 74773
rect 29729 74745 29763 74773
rect 29791 74745 32619 74773
rect 32647 74745 32681 74773
rect 32709 74745 47979 74773
rect 48007 74745 48041 74773
rect 48069 74745 63339 74773
rect 63367 74745 63401 74773
rect 63429 74745 78699 74773
rect 78727 74745 78761 74773
rect 78789 74745 94059 74773
rect 94087 74745 94121 74773
rect 94149 74745 109419 74773
rect 109447 74745 109481 74773
rect 109509 74745 124779 74773
rect 124807 74745 124841 74773
rect 124869 74745 140139 74773
rect 140167 74745 140201 74773
rect 140229 74745 155499 74773
rect 155527 74745 155561 74773
rect 155589 74745 170859 74773
rect 170887 74745 170921 74773
rect 170949 74745 186219 74773
rect 186247 74745 186281 74773
rect 186309 74745 201579 74773
rect 201607 74745 201641 74773
rect 201669 74745 216939 74773
rect 216967 74745 217001 74773
rect 217029 74745 232299 74773
rect 232327 74745 232361 74773
rect 232389 74745 247659 74773
rect 247687 74745 247721 74773
rect 247749 74745 254577 74773
rect 254605 74745 254639 74773
rect 254667 74745 254701 74773
rect 254729 74745 254763 74773
rect 254791 74745 263577 74773
rect 263605 74745 263639 74773
rect 263667 74745 263701 74773
rect 263729 74745 263763 74773
rect 263791 74745 272577 74773
rect 272605 74745 272639 74773
rect 272667 74745 272701 74773
rect 272729 74745 272763 74773
rect 272791 74745 281577 74773
rect 281605 74745 281639 74773
rect 281667 74745 281701 74773
rect 281729 74745 281763 74773
rect 281791 74745 290577 74773
rect 290605 74745 290639 74773
rect 290667 74745 290701 74773
rect 290729 74745 290763 74773
rect 290791 74745 299256 74773
rect 299284 74745 299318 74773
rect 299346 74745 299380 74773
rect 299408 74745 299442 74773
rect 299470 74745 299998 74773
rect -6 74697 299998 74745
rect -6 68959 299998 69007
rect -6 68931 42 68959
rect 70 68931 104 68959
rect 132 68931 166 68959
rect 194 68931 228 68959
rect 256 68931 4437 68959
rect 4465 68931 4499 68959
rect 4527 68931 4561 68959
rect 4589 68931 4623 68959
rect 4651 68931 13437 68959
rect 13465 68931 13499 68959
rect 13527 68931 13561 68959
rect 13589 68931 13623 68959
rect 13651 68931 22437 68959
rect 22465 68931 22499 68959
rect 22527 68931 22561 68959
rect 22589 68931 22623 68959
rect 22651 68931 24939 68959
rect 24967 68931 25001 68959
rect 25029 68931 31437 68959
rect 31465 68931 31499 68959
rect 31527 68931 31561 68959
rect 31589 68931 31623 68959
rect 31651 68931 40299 68959
rect 40327 68931 40361 68959
rect 40389 68931 55659 68959
rect 55687 68931 55721 68959
rect 55749 68931 71019 68959
rect 71047 68931 71081 68959
rect 71109 68931 86379 68959
rect 86407 68931 86441 68959
rect 86469 68931 101739 68959
rect 101767 68931 101801 68959
rect 101829 68931 117099 68959
rect 117127 68931 117161 68959
rect 117189 68931 132459 68959
rect 132487 68931 132521 68959
rect 132549 68931 147819 68959
rect 147847 68931 147881 68959
rect 147909 68931 163179 68959
rect 163207 68931 163241 68959
rect 163269 68931 178539 68959
rect 178567 68931 178601 68959
rect 178629 68931 193899 68959
rect 193927 68931 193961 68959
rect 193989 68931 209259 68959
rect 209287 68931 209321 68959
rect 209349 68931 224619 68959
rect 224647 68931 224681 68959
rect 224709 68931 239979 68959
rect 240007 68931 240041 68959
rect 240069 68931 256437 68959
rect 256465 68931 256499 68959
rect 256527 68931 256561 68959
rect 256589 68931 256623 68959
rect 256651 68931 265437 68959
rect 265465 68931 265499 68959
rect 265527 68931 265561 68959
rect 265589 68931 265623 68959
rect 265651 68931 274437 68959
rect 274465 68931 274499 68959
rect 274527 68931 274561 68959
rect 274589 68931 274623 68959
rect 274651 68931 283437 68959
rect 283465 68931 283499 68959
rect 283527 68931 283561 68959
rect 283589 68931 283623 68959
rect 283651 68931 292437 68959
rect 292465 68931 292499 68959
rect 292527 68931 292561 68959
rect 292589 68931 292623 68959
rect 292651 68931 299736 68959
rect 299764 68931 299798 68959
rect 299826 68931 299860 68959
rect 299888 68931 299922 68959
rect 299950 68931 299998 68959
rect -6 68897 299998 68931
rect -6 68869 42 68897
rect 70 68869 104 68897
rect 132 68869 166 68897
rect 194 68869 228 68897
rect 256 68869 4437 68897
rect 4465 68869 4499 68897
rect 4527 68869 4561 68897
rect 4589 68869 4623 68897
rect 4651 68869 13437 68897
rect 13465 68869 13499 68897
rect 13527 68869 13561 68897
rect 13589 68869 13623 68897
rect 13651 68869 22437 68897
rect 22465 68869 22499 68897
rect 22527 68869 22561 68897
rect 22589 68869 22623 68897
rect 22651 68869 24939 68897
rect 24967 68869 25001 68897
rect 25029 68869 31437 68897
rect 31465 68869 31499 68897
rect 31527 68869 31561 68897
rect 31589 68869 31623 68897
rect 31651 68869 40299 68897
rect 40327 68869 40361 68897
rect 40389 68869 55659 68897
rect 55687 68869 55721 68897
rect 55749 68869 71019 68897
rect 71047 68869 71081 68897
rect 71109 68869 86379 68897
rect 86407 68869 86441 68897
rect 86469 68869 101739 68897
rect 101767 68869 101801 68897
rect 101829 68869 117099 68897
rect 117127 68869 117161 68897
rect 117189 68869 132459 68897
rect 132487 68869 132521 68897
rect 132549 68869 147819 68897
rect 147847 68869 147881 68897
rect 147909 68869 163179 68897
rect 163207 68869 163241 68897
rect 163269 68869 178539 68897
rect 178567 68869 178601 68897
rect 178629 68869 193899 68897
rect 193927 68869 193961 68897
rect 193989 68869 209259 68897
rect 209287 68869 209321 68897
rect 209349 68869 224619 68897
rect 224647 68869 224681 68897
rect 224709 68869 239979 68897
rect 240007 68869 240041 68897
rect 240069 68869 256437 68897
rect 256465 68869 256499 68897
rect 256527 68869 256561 68897
rect 256589 68869 256623 68897
rect 256651 68869 265437 68897
rect 265465 68869 265499 68897
rect 265527 68869 265561 68897
rect 265589 68869 265623 68897
rect 265651 68869 274437 68897
rect 274465 68869 274499 68897
rect 274527 68869 274561 68897
rect 274589 68869 274623 68897
rect 274651 68869 283437 68897
rect 283465 68869 283499 68897
rect 283527 68869 283561 68897
rect 283589 68869 283623 68897
rect 283651 68869 292437 68897
rect 292465 68869 292499 68897
rect 292527 68869 292561 68897
rect 292589 68869 292623 68897
rect 292651 68869 299736 68897
rect 299764 68869 299798 68897
rect 299826 68869 299860 68897
rect 299888 68869 299922 68897
rect 299950 68869 299998 68897
rect -6 68835 299998 68869
rect -6 68807 42 68835
rect 70 68807 104 68835
rect 132 68807 166 68835
rect 194 68807 228 68835
rect 256 68807 4437 68835
rect 4465 68807 4499 68835
rect 4527 68807 4561 68835
rect 4589 68807 4623 68835
rect 4651 68807 13437 68835
rect 13465 68807 13499 68835
rect 13527 68807 13561 68835
rect 13589 68807 13623 68835
rect 13651 68807 22437 68835
rect 22465 68807 22499 68835
rect 22527 68807 22561 68835
rect 22589 68807 22623 68835
rect 22651 68807 24939 68835
rect 24967 68807 25001 68835
rect 25029 68807 31437 68835
rect 31465 68807 31499 68835
rect 31527 68807 31561 68835
rect 31589 68807 31623 68835
rect 31651 68807 40299 68835
rect 40327 68807 40361 68835
rect 40389 68807 55659 68835
rect 55687 68807 55721 68835
rect 55749 68807 71019 68835
rect 71047 68807 71081 68835
rect 71109 68807 86379 68835
rect 86407 68807 86441 68835
rect 86469 68807 101739 68835
rect 101767 68807 101801 68835
rect 101829 68807 117099 68835
rect 117127 68807 117161 68835
rect 117189 68807 132459 68835
rect 132487 68807 132521 68835
rect 132549 68807 147819 68835
rect 147847 68807 147881 68835
rect 147909 68807 163179 68835
rect 163207 68807 163241 68835
rect 163269 68807 178539 68835
rect 178567 68807 178601 68835
rect 178629 68807 193899 68835
rect 193927 68807 193961 68835
rect 193989 68807 209259 68835
rect 209287 68807 209321 68835
rect 209349 68807 224619 68835
rect 224647 68807 224681 68835
rect 224709 68807 239979 68835
rect 240007 68807 240041 68835
rect 240069 68807 256437 68835
rect 256465 68807 256499 68835
rect 256527 68807 256561 68835
rect 256589 68807 256623 68835
rect 256651 68807 265437 68835
rect 265465 68807 265499 68835
rect 265527 68807 265561 68835
rect 265589 68807 265623 68835
rect 265651 68807 274437 68835
rect 274465 68807 274499 68835
rect 274527 68807 274561 68835
rect 274589 68807 274623 68835
rect 274651 68807 283437 68835
rect 283465 68807 283499 68835
rect 283527 68807 283561 68835
rect 283589 68807 283623 68835
rect 283651 68807 292437 68835
rect 292465 68807 292499 68835
rect 292527 68807 292561 68835
rect 292589 68807 292623 68835
rect 292651 68807 299736 68835
rect 299764 68807 299798 68835
rect 299826 68807 299860 68835
rect 299888 68807 299922 68835
rect 299950 68807 299998 68835
rect -6 68773 299998 68807
rect -6 68745 42 68773
rect 70 68745 104 68773
rect 132 68745 166 68773
rect 194 68745 228 68773
rect 256 68745 4437 68773
rect 4465 68745 4499 68773
rect 4527 68745 4561 68773
rect 4589 68745 4623 68773
rect 4651 68745 13437 68773
rect 13465 68745 13499 68773
rect 13527 68745 13561 68773
rect 13589 68745 13623 68773
rect 13651 68745 22437 68773
rect 22465 68745 22499 68773
rect 22527 68745 22561 68773
rect 22589 68745 22623 68773
rect 22651 68745 24939 68773
rect 24967 68745 25001 68773
rect 25029 68745 31437 68773
rect 31465 68745 31499 68773
rect 31527 68745 31561 68773
rect 31589 68745 31623 68773
rect 31651 68745 40299 68773
rect 40327 68745 40361 68773
rect 40389 68745 55659 68773
rect 55687 68745 55721 68773
rect 55749 68745 71019 68773
rect 71047 68745 71081 68773
rect 71109 68745 86379 68773
rect 86407 68745 86441 68773
rect 86469 68745 101739 68773
rect 101767 68745 101801 68773
rect 101829 68745 117099 68773
rect 117127 68745 117161 68773
rect 117189 68745 132459 68773
rect 132487 68745 132521 68773
rect 132549 68745 147819 68773
rect 147847 68745 147881 68773
rect 147909 68745 163179 68773
rect 163207 68745 163241 68773
rect 163269 68745 178539 68773
rect 178567 68745 178601 68773
rect 178629 68745 193899 68773
rect 193927 68745 193961 68773
rect 193989 68745 209259 68773
rect 209287 68745 209321 68773
rect 209349 68745 224619 68773
rect 224647 68745 224681 68773
rect 224709 68745 239979 68773
rect 240007 68745 240041 68773
rect 240069 68745 256437 68773
rect 256465 68745 256499 68773
rect 256527 68745 256561 68773
rect 256589 68745 256623 68773
rect 256651 68745 265437 68773
rect 265465 68745 265499 68773
rect 265527 68745 265561 68773
rect 265589 68745 265623 68773
rect 265651 68745 274437 68773
rect 274465 68745 274499 68773
rect 274527 68745 274561 68773
rect 274589 68745 274623 68773
rect 274651 68745 283437 68773
rect 283465 68745 283499 68773
rect 283527 68745 283561 68773
rect 283589 68745 283623 68773
rect 283651 68745 292437 68773
rect 292465 68745 292499 68773
rect 292527 68745 292561 68773
rect 292589 68745 292623 68773
rect 292651 68745 299736 68773
rect 299764 68745 299798 68773
rect 299826 68745 299860 68773
rect 299888 68745 299922 68773
rect 299950 68745 299998 68773
rect -6 68697 299998 68745
rect -6 65959 299998 66007
rect -6 65931 522 65959
rect 550 65931 584 65959
rect 612 65931 646 65959
rect 674 65931 708 65959
rect 736 65931 2577 65959
rect 2605 65931 2639 65959
rect 2667 65931 2701 65959
rect 2729 65931 2763 65959
rect 2791 65931 11577 65959
rect 11605 65931 11639 65959
rect 11667 65931 11701 65959
rect 11729 65931 11763 65959
rect 11791 65931 17259 65959
rect 17287 65931 17321 65959
rect 17349 65931 20577 65959
rect 20605 65931 20639 65959
rect 20667 65931 20701 65959
rect 20729 65931 20763 65959
rect 20791 65931 29577 65959
rect 29605 65931 29639 65959
rect 29667 65931 29701 65959
rect 29729 65931 29763 65959
rect 29791 65931 32619 65959
rect 32647 65931 32681 65959
rect 32709 65931 47979 65959
rect 48007 65931 48041 65959
rect 48069 65931 63339 65959
rect 63367 65931 63401 65959
rect 63429 65931 78699 65959
rect 78727 65931 78761 65959
rect 78789 65931 94059 65959
rect 94087 65931 94121 65959
rect 94149 65931 109419 65959
rect 109447 65931 109481 65959
rect 109509 65931 124779 65959
rect 124807 65931 124841 65959
rect 124869 65931 140139 65959
rect 140167 65931 140201 65959
rect 140229 65931 155499 65959
rect 155527 65931 155561 65959
rect 155589 65931 170859 65959
rect 170887 65931 170921 65959
rect 170949 65931 186219 65959
rect 186247 65931 186281 65959
rect 186309 65931 201579 65959
rect 201607 65931 201641 65959
rect 201669 65931 216939 65959
rect 216967 65931 217001 65959
rect 217029 65931 232299 65959
rect 232327 65931 232361 65959
rect 232389 65931 247659 65959
rect 247687 65931 247721 65959
rect 247749 65931 254577 65959
rect 254605 65931 254639 65959
rect 254667 65931 254701 65959
rect 254729 65931 254763 65959
rect 254791 65931 263577 65959
rect 263605 65931 263639 65959
rect 263667 65931 263701 65959
rect 263729 65931 263763 65959
rect 263791 65931 272577 65959
rect 272605 65931 272639 65959
rect 272667 65931 272701 65959
rect 272729 65931 272763 65959
rect 272791 65931 281577 65959
rect 281605 65931 281639 65959
rect 281667 65931 281701 65959
rect 281729 65931 281763 65959
rect 281791 65931 290577 65959
rect 290605 65931 290639 65959
rect 290667 65931 290701 65959
rect 290729 65931 290763 65959
rect 290791 65931 299256 65959
rect 299284 65931 299318 65959
rect 299346 65931 299380 65959
rect 299408 65931 299442 65959
rect 299470 65931 299998 65959
rect -6 65897 299998 65931
rect -6 65869 522 65897
rect 550 65869 584 65897
rect 612 65869 646 65897
rect 674 65869 708 65897
rect 736 65869 2577 65897
rect 2605 65869 2639 65897
rect 2667 65869 2701 65897
rect 2729 65869 2763 65897
rect 2791 65869 11577 65897
rect 11605 65869 11639 65897
rect 11667 65869 11701 65897
rect 11729 65869 11763 65897
rect 11791 65869 17259 65897
rect 17287 65869 17321 65897
rect 17349 65869 20577 65897
rect 20605 65869 20639 65897
rect 20667 65869 20701 65897
rect 20729 65869 20763 65897
rect 20791 65869 29577 65897
rect 29605 65869 29639 65897
rect 29667 65869 29701 65897
rect 29729 65869 29763 65897
rect 29791 65869 32619 65897
rect 32647 65869 32681 65897
rect 32709 65869 47979 65897
rect 48007 65869 48041 65897
rect 48069 65869 63339 65897
rect 63367 65869 63401 65897
rect 63429 65869 78699 65897
rect 78727 65869 78761 65897
rect 78789 65869 94059 65897
rect 94087 65869 94121 65897
rect 94149 65869 109419 65897
rect 109447 65869 109481 65897
rect 109509 65869 124779 65897
rect 124807 65869 124841 65897
rect 124869 65869 140139 65897
rect 140167 65869 140201 65897
rect 140229 65869 155499 65897
rect 155527 65869 155561 65897
rect 155589 65869 170859 65897
rect 170887 65869 170921 65897
rect 170949 65869 186219 65897
rect 186247 65869 186281 65897
rect 186309 65869 201579 65897
rect 201607 65869 201641 65897
rect 201669 65869 216939 65897
rect 216967 65869 217001 65897
rect 217029 65869 232299 65897
rect 232327 65869 232361 65897
rect 232389 65869 247659 65897
rect 247687 65869 247721 65897
rect 247749 65869 254577 65897
rect 254605 65869 254639 65897
rect 254667 65869 254701 65897
rect 254729 65869 254763 65897
rect 254791 65869 263577 65897
rect 263605 65869 263639 65897
rect 263667 65869 263701 65897
rect 263729 65869 263763 65897
rect 263791 65869 272577 65897
rect 272605 65869 272639 65897
rect 272667 65869 272701 65897
rect 272729 65869 272763 65897
rect 272791 65869 281577 65897
rect 281605 65869 281639 65897
rect 281667 65869 281701 65897
rect 281729 65869 281763 65897
rect 281791 65869 290577 65897
rect 290605 65869 290639 65897
rect 290667 65869 290701 65897
rect 290729 65869 290763 65897
rect 290791 65869 299256 65897
rect 299284 65869 299318 65897
rect 299346 65869 299380 65897
rect 299408 65869 299442 65897
rect 299470 65869 299998 65897
rect -6 65835 299998 65869
rect -6 65807 522 65835
rect 550 65807 584 65835
rect 612 65807 646 65835
rect 674 65807 708 65835
rect 736 65807 2577 65835
rect 2605 65807 2639 65835
rect 2667 65807 2701 65835
rect 2729 65807 2763 65835
rect 2791 65807 11577 65835
rect 11605 65807 11639 65835
rect 11667 65807 11701 65835
rect 11729 65807 11763 65835
rect 11791 65807 17259 65835
rect 17287 65807 17321 65835
rect 17349 65807 20577 65835
rect 20605 65807 20639 65835
rect 20667 65807 20701 65835
rect 20729 65807 20763 65835
rect 20791 65807 29577 65835
rect 29605 65807 29639 65835
rect 29667 65807 29701 65835
rect 29729 65807 29763 65835
rect 29791 65807 32619 65835
rect 32647 65807 32681 65835
rect 32709 65807 47979 65835
rect 48007 65807 48041 65835
rect 48069 65807 63339 65835
rect 63367 65807 63401 65835
rect 63429 65807 78699 65835
rect 78727 65807 78761 65835
rect 78789 65807 94059 65835
rect 94087 65807 94121 65835
rect 94149 65807 109419 65835
rect 109447 65807 109481 65835
rect 109509 65807 124779 65835
rect 124807 65807 124841 65835
rect 124869 65807 140139 65835
rect 140167 65807 140201 65835
rect 140229 65807 155499 65835
rect 155527 65807 155561 65835
rect 155589 65807 170859 65835
rect 170887 65807 170921 65835
rect 170949 65807 186219 65835
rect 186247 65807 186281 65835
rect 186309 65807 201579 65835
rect 201607 65807 201641 65835
rect 201669 65807 216939 65835
rect 216967 65807 217001 65835
rect 217029 65807 232299 65835
rect 232327 65807 232361 65835
rect 232389 65807 247659 65835
rect 247687 65807 247721 65835
rect 247749 65807 254577 65835
rect 254605 65807 254639 65835
rect 254667 65807 254701 65835
rect 254729 65807 254763 65835
rect 254791 65807 263577 65835
rect 263605 65807 263639 65835
rect 263667 65807 263701 65835
rect 263729 65807 263763 65835
rect 263791 65807 272577 65835
rect 272605 65807 272639 65835
rect 272667 65807 272701 65835
rect 272729 65807 272763 65835
rect 272791 65807 281577 65835
rect 281605 65807 281639 65835
rect 281667 65807 281701 65835
rect 281729 65807 281763 65835
rect 281791 65807 290577 65835
rect 290605 65807 290639 65835
rect 290667 65807 290701 65835
rect 290729 65807 290763 65835
rect 290791 65807 299256 65835
rect 299284 65807 299318 65835
rect 299346 65807 299380 65835
rect 299408 65807 299442 65835
rect 299470 65807 299998 65835
rect -6 65773 299998 65807
rect -6 65745 522 65773
rect 550 65745 584 65773
rect 612 65745 646 65773
rect 674 65745 708 65773
rect 736 65745 2577 65773
rect 2605 65745 2639 65773
rect 2667 65745 2701 65773
rect 2729 65745 2763 65773
rect 2791 65745 11577 65773
rect 11605 65745 11639 65773
rect 11667 65745 11701 65773
rect 11729 65745 11763 65773
rect 11791 65745 17259 65773
rect 17287 65745 17321 65773
rect 17349 65745 20577 65773
rect 20605 65745 20639 65773
rect 20667 65745 20701 65773
rect 20729 65745 20763 65773
rect 20791 65745 29577 65773
rect 29605 65745 29639 65773
rect 29667 65745 29701 65773
rect 29729 65745 29763 65773
rect 29791 65745 32619 65773
rect 32647 65745 32681 65773
rect 32709 65745 47979 65773
rect 48007 65745 48041 65773
rect 48069 65745 63339 65773
rect 63367 65745 63401 65773
rect 63429 65745 78699 65773
rect 78727 65745 78761 65773
rect 78789 65745 94059 65773
rect 94087 65745 94121 65773
rect 94149 65745 109419 65773
rect 109447 65745 109481 65773
rect 109509 65745 124779 65773
rect 124807 65745 124841 65773
rect 124869 65745 140139 65773
rect 140167 65745 140201 65773
rect 140229 65745 155499 65773
rect 155527 65745 155561 65773
rect 155589 65745 170859 65773
rect 170887 65745 170921 65773
rect 170949 65745 186219 65773
rect 186247 65745 186281 65773
rect 186309 65745 201579 65773
rect 201607 65745 201641 65773
rect 201669 65745 216939 65773
rect 216967 65745 217001 65773
rect 217029 65745 232299 65773
rect 232327 65745 232361 65773
rect 232389 65745 247659 65773
rect 247687 65745 247721 65773
rect 247749 65745 254577 65773
rect 254605 65745 254639 65773
rect 254667 65745 254701 65773
rect 254729 65745 254763 65773
rect 254791 65745 263577 65773
rect 263605 65745 263639 65773
rect 263667 65745 263701 65773
rect 263729 65745 263763 65773
rect 263791 65745 272577 65773
rect 272605 65745 272639 65773
rect 272667 65745 272701 65773
rect 272729 65745 272763 65773
rect 272791 65745 281577 65773
rect 281605 65745 281639 65773
rect 281667 65745 281701 65773
rect 281729 65745 281763 65773
rect 281791 65745 290577 65773
rect 290605 65745 290639 65773
rect 290667 65745 290701 65773
rect 290729 65745 290763 65773
rect 290791 65745 299256 65773
rect 299284 65745 299318 65773
rect 299346 65745 299380 65773
rect 299408 65745 299442 65773
rect 299470 65745 299998 65773
rect -6 65697 299998 65745
rect -6 59959 299998 60007
rect -6 59931 42 59959
rect 70 59931 104 59959
rect 132 59931 166 59959
rect 194 59931 228 59959
rect 256 59931 4437 59959
rect 4465 59931 4499 59959
rect 4527 59931 4561 59959
rect 4589 59931 4623 59959
rect 4651 59931 13437 59959
rect 13465 59931 13499 59959
rect 13527 59931 13561 59959
rect 13589 59931 13623 59959
rect 13651 59931 22437 59959
rect 22465 59931 22499 59959
rect 22527 59931 22561 59959
rect 22589 59931 22623 59959
rect 22651 59931 24939 59959
rect 24967 59931 25001 59959
rect 25029 59931 31437 59959
rect 31465 59931 31499 59959
rect 31527 59931 31561 59959
rect 31589 59931 31623 59959
rect 31651 59931 40299 59959
rect 40327 59931 40361 59959
rect 40389 59931 55659 59959
rect 55687 59931 55721 59959
rect 55749 59931 71019 59959
rect 71047 59931 71081 59959
rect 71109 59931 86379 59959
rect 86407 59931 86441 59959
rect 86469 59931 101739 59959
rect 101767 59931 101801 59959
rect 101829 59931 117099 59959
rect 117127 59931 117161 59959
rect 117189 59931 132459 59959
rect 132487 59931 132521 59959
rect 132549 59931 147819 59959
rect 147847 59931 147881 59959
rect 147909 59931 163179 59959
rect 163207 59931 163241 59959
rect 163269 59931 178539 59959
rect 178567 59931 178601 59959
rect 178629 59931 193899 59959
rect 193927 59931 193961 59959
rect 193989 59931 209259 59959
rect 209287 59931 209321 59959
rect 209349 59931 224619 59959
rect 224647 59931 224681 59959
rect 224709 59931 239979 59959
rect 240007 59931 240041 59959
rect 240069 59931 256437 59959
rect 256465 59931 256499 59959
rect 256527 59931 256561 59959
rect 256589 59931 256623 59959
rect 256651 59931 265437 59959
rect 265465 59931 265499 59959
rect 265527 59931 265561 59959
rect 265589 59931 265623 59959
rect 265651 59931 274437 59959
rect 274465 59931 274499 59959
rect 274527 59931 274561 59959
rect 274589 59931 274623 59959
rect 274651 59931 283437 59959
rect 283465 59931 283499 59959
rect 283527 59931 283561 59959
rect 283589 59931 283623 59959
rect 283651 59931 292437 59959
rect 292465 59931 292499 59959
rect 292527 59931 292561 59959
rect 292589 59931 292623 59959
rect 292651 59931 299736 59959
rect 299764 59931 299798 59959
rect 299826 59931 299860 59959
rect 299888 59931 299922 59959
rect 299950 59931 299998 59959
rect -6 59897 299998 59931
rect -6 59869 42 59897
rect 70 59869 104 59897
rect 132 59869 166 59897
rect 194 59869 228 59897
rect 256 59869 4437 59897
rect 4465 59869 4499 59897
rect 4527 59869 4561 59897
rect 4589 59869 4623 59897
rect 4651 59869 13437 59897
rect 13465 59869 13499 59897
rect 13527 59869 13561 59897
rect 13589 59869 13623 59897
rect 13651 59869 22437 59897
rect 22465 59869 22499 59897
rect 22527 59869 22561 59897
rect 22589 59869 22623 59897
rect 22651 59869 24939 59897
rect 24967 59869 25001 59897
rect 25029 59869 31437 59897
rect 31465 59869 31499 59897
rect 31527 59869 31561 59897
rect 31589 59869 31623 59897
rect 31651 59869 40299 59897
rect 40327 59869 40361 59897
rect 40389 59869 55659 59897
rect 55687 59869 55721 59897
rect 55749 59869 71019 59897
rect 71047 59869 71081 59897
rect 71109 59869 86379 59897
rect 86407 59869 86441 59897
rect 86469 59869 101739 59897
rect 101767 59869 101801 59897
rect 101829 59869 117099 59897
rect 117127 59869 117161 59897
rect 117189 59869 132459 59897
rect 132487 59869 132521 59897
rect 132549 59869 147819 59897
rect 147847 59869 147881 59897
rect 147909 59869 163179 59897
rect 163207 59869 163241 59897
rect 163269 59869 178539 59897
rect 178567 59869 178601 59897
rect 178629 59869 193899 59897
rect 193927 59869 193961 59897
rect 193989 59869 209259 59897
rect 209287 59869 209321 59897
rect 209349 59869 224619 59897
rect 224647 59869 224681 59897
rect 224709 59869 239979 59897
rect 240007 59869 240041 59897
rect 240069 59869 256437 59897
rect 256465 59869 256499 59897
rect 256527 59869 256561 59897
rect 256589 59869 256623 59897
rect 256651 59869 265437 59897
rect 265465 59869 265499 59897
rect 265527 59869 265561 59897
rect 265589 59869 265623 59897
rect 265651 59869 274437 59897
rect 274465 59869 274499 59897
rect 274527 59869 274561 59897
rect 274589 59869 274623 59897
rect 274651 59869 283437 59897
rect 283465 59869 283499 59897
rect 283527 59869 283561 59897
rect 283589 59869 283623 59897
rect 283651 59869 292437 59897
rect 292465 59869 292499 59897
rect 292527 59869 292561 59897
rect 292589 59869 292623 59897
rect 292651 59869 299736 59897
rect 299764 59869 299798 59897
rect 299826 59869 299860 59897
rect 299888 59869 299922 59897
rect 299950 59869 299998 59897
rect -6 59835 299998 59869
rect -6 59807 42 59835
rect 70 59807 104 59835
rect 132 59807 166 59835
rect 194 59807 228 59835
rect 256 59807 4437 59835
rect 4465 59807 4499 59835
rect 4527 59807 4561 59835
rect 4589 59807 4623 59835
rect 4651 59807 13437 59835
rect 13465 59807 13499 59835
rect 13527 59807 13561 59835
rect 13589 59807 13623 59835
rect 13651 59807 22437 59835
rect 22465 59807 22499 59835
rect 22527 59807 22561 59835
rect 22589 59807 22623 59835
rect 22651 59807 24939 59835
rect 24967 59807 25001 59835
rect 25029 59807 31437 59835
rect 31465 59807 31499 59835
rect 31527 59807 31561 59835
rect 31589 59807 31623 59835
rect 31651 59807 40299 59835
rect 40327 59807 40361 59835
rect 40389 59807 55659 59835
rect 55687 59807 55721 59835
rect 55749 59807 71019 59835
rect 71047 59807 71081 59835
rect 71109 59807 86379 59835
rect 86407 59807 86441 59835
rect 86469 59807 101739 59835
rect 101767 59807 101801 59835
rect 101829 59807 117099 59835
rect 117127 59807 117161 59835
rect 117189 59807 132459 59835
rect 132487 59807 132521 59835
rect 132549 59807 147819 59835
rect 147847 59807 147881 59835
rect 147909 59807 163179 59835
rect 163207 59807 163241 59835
rect 163269 59807 178539 59835
rect 178567 59807 178601 59835
rect 178629 59807 193899 59835
rect 193927 59807 193961 59835
rect 193989 59807 209259 59835
rect 209287 59807 209321 59835
rect 209349 59807 224619 59835
rect 224647 59807 224681 59835
rect 224709 59807 239979 59835
rect 240007 59807 240041 59835
rect 240069 59807 256437 59835
rect 256465 59807 256499 59835
rect 256527 59807 256561 59835
rect 256589 59807 256623 59835
rect 256651 59807 265437 59835
rect 265465 59807 265499 59835
rect 265527 59807 265561 59835
rect 265589 59807 265623 59835
rect 265651 59807 274437 59835
rect 274465 59807 274499 59835
rect 274527 59807 274561 59835
rect 274589 59807 274623 59835
rect 274651 59807 283437 59835
rect 283465 59807 283499 59835
rect 283527 59807 283561 59835
rect 283589 59807 283623 59835
rect 283651 59807 292437 59835
rect 292465 59807 292499 59835
rect 292527 59807 292561 59835
rect 292589 59807 292623 59835
rect 292651 59807 299736 59835
rect 299764 59807 299798 59835
rect 299826 59807 299860 59835
rect 299888 59807 299922 59835
rect 299950 59807 299998 59835
rect -6 59773 299998 59807
rect -6 59745 42 59773
rect 70 59745 104 59773
rect 132 59745 166 59773
rect 194 59745 228 59773
rect 256 59745 4437 59773
rect 4465 59745 4499 59773
rect 4527 59745 4561 59773
rect 4589 59745 4623 59773
rect 4651 59745 13437 59773
rect 13465 59745 13499 59773
rect 13527 59745 13561 59773
rect 13589 59745 13623 59773
rect 13651 59745 22437 59773
rect 22465 59745 22499 59773
rect 22527 59745 22561 59773
rect 22589 59745 22623 59773
rect 22651 59745 24939 59773
rect 24967 59745 25001 59773
rect 25029 59745 31437 59773
rect 31465 59745 31499 59773
rect 31527 59745 31561 59773
rect 31589 59745 31623 59773
rect 31651 59745 40299 59773
rect 40327 59745 40361 59773
rect 40389 59745 55659 59773
rect 55687 59745 55721 59773
rect 55749 59745 71019 59773
rect 71047 59745 71081 59773
rect 71109 59745 86379 59773
rect 86407 59745 86441 59773
rect 86469 59745 101739 59773
rect 101767 59745 101801 59773
rect 101829 59745 117099 59773
rect 117127 59745 117161 59773
rect 117189 59745 132459 59773
rect 132487 59745 132521 59773
rect 132549 59745 147819 59773
rect 147847 59745 147881 59773
rect 147909 59745 163179 59773
rect 163207 59745 163241 59773
rect 163269 59745 178539 59773
rect 178567 59745 178601 59773
rect 178629 59745 193899 59773
rect 193927 59745 193961 59773
rect 193989 59745 209259 59773
rect 209287 59745 209321 59773
rect 209349 59745 224619 59773
rect 224647 59745 224681 59773
rect 224709 59745 239979 59773
rect 240007 59745 240041 59773
rect 240069 59745 256437 59773
rect 256465 59745 256499 59773
rect 256527 59745 256561 59773
rect 256589 59745 256623 59773
rect 256651 59745 265437 59773
rect 265465 59745 265499 59773
rect 265527 59745 265561 59773
rect 265589 59745 265623 59773
rect 265651 59745 274437 59773
rect 274465 59745 274499 59773
rect 274527 59745 274561 59773
rect 274589 59745 274623 59773
rect 274651 59745 283437 59773
rect 283465 59745 283499 59773
rect 283527 59745 283561 59773
rect 283589 59745 283623 59773
rect 283651 59745 292437 59773
rect 292465 59745 292499 59773
rect 292527 59745 292561 59773
rect 292589 59745 292623 59773
rect 292651 59745 299736 59773
rect 299764 59745 299798 59773
rect 299826 59745 299860 59773
rect 299888 59745 299922 59773
rect 299950 59745 299998 59773
rect -6 59697 299998 59745
rect -6 56959 299998 57007
rect -6 56931 522 56959
rect 550 56931 584 56959
rect 612 56931 646 56959
rect 674 56931 708 56959
rect 736 56931 2577 56959
rect 2605 56931 2639 56959
rect 2667 56931 2701 56959
rect 2729 56931 2763 56959
rect 2791 56931 11577 56959
rect 11605 56931 11639 56959
rect 11667 56931 11701 56959
rect 11729 56931 11763 56959
rect 11791 56931 17259 56959
rect 17287 56931 17321 56959
rect 17349 56931 20577 56959
rect 20605 56931 20639 56959
rect 20667 56931 20701 56959
rect 20729 56931 20763 56959
rect 20791 56931 29577 56959
rect 29605 56931 29639 56959
rect 29667 56931 29701 56959
rect 29729 56931 29763 56959
rect 29791 56931 32619 56959
rect 32647 56931 32681 56959
rect 32709 56931 47979 56959
rect 48007 56931 48041 56959
rect 48069 56931 63339 56959
rect 63367 56931 63401 56959
rect 63429 56931 78699 56959
rect 78727 56931 78761 56959
rect 78789 56931 94059 56959
rect 94087 56931 94121 56959
rect 94149 56931 109419 56959
rect 109447 56931 109481 56959
rect 109509 56931 124779 56959
rect 124807 56931 124841 56959
rect 124869 56931 140139 56959
rect 140167 56931 140201 56959
rect 140229 56931 155499 56959
rect 155527 56931 155561 56959
rect 155589 56931 170859 56959
rect 170887 56931 170921 56959
rect 170949 56931 186219 56959
rect 186247 56931 186281 56959
rect 186309 56931 201579 56959
rect 201607 56931 201641 56959
rect 201669 56931 216939 56959
rect 216967 56931 217001 56959
rect 217029 56931 232299 56959
rect 232327 56931 232361 56959
rect 232389 56931 247659 56959
rect 247687 56931 247721 56959
rect 247749 56931 254577 56959
rect 254605 56931 254639 56959
rect 254667 56931 254701 56959
rect 254729 56931 254763 56959
rect 254791 56931 263577 56959
rect 263605 56931 263639 56959
rect 263667 56931 263701 56959
rect 263729 56931 263763 56959
rect 263791 56931 272577 56959
rect 272605 56931 272639 56959
rect 272667 56931 272701 56959
rect 272729 56931 272763 56959
rect 272791 56931 281577 56959
rect 281605 56931 281639 56959
rect 281667 56931 281701 56959
rect 281729 56931 281763 56959
rect 281791 56931 290577 56959
rect 290605 56931 290639 56959
rect 290667 56931 290701 56959
rect 290729 56931 290763 56959
rect 290791 56931 299256 56959
rect 299284 56931 299318 56959
rect 299346 56931 299380 56959
rect 299408 56931 299442 56959
rect 299470 56931 299998 56959
rect -6 56897 299998 56931
rect -6 56869 522 56897
rect 550 56869 584 56897
rect 612 56869 646 56897
rect 674 56869 708 56897
rect 736 56869 2577 56897
rect 2605 56869 2639 56897
rect 2667 56869 2701 56897
rect 2729 56869 2763 56897
rect 2791 56869 11577 56897
rect 11605 56869 11639 56897
rect 11667 56869 11701 56897
rect 11729 56869 11763 56897
rect 11791 56869 17259 56897
rect 17287 56869 17321 56897
rect 17349 56869 20577 56897
rect 20605 56869 20639 56897
rect 20667 56869 20701 56897
rect 20729 56869 20763 56897
rect 20791 56869 29577 56897
rect 29605 56869 29639 56897
rect 29667 56869 29701 56897
rect 29729 56869 29763 56897
rect 29791 56869 32619 56897
rect 32647 56869 32681 56897
rect 32709 56869 47979 56897
rect 48007 56869 48041 56897
rect 48069 56869 63339 56897
rect 63367 56869 63401 56897
rect 63429 56869 78699 56897
rect 78727 56869 78761 56897
rect 78789 56869 94059 56897
rect 94087 56869 94121 56897
rect 94149 56869 109419 56897
rect 109447 56869 109481 56897
rect 109509 56869 124779 56897
rect 124807 56869 124841 56897
rect 124869 56869 140139 56897
rect 140167 56869 140201 56897
rect 140229 56869 155499 56897
rect 155527 56869 155561 56897
rect 155589 56869 170859 56897
rect 170887 56869 170921 56897
rect 170949 56869 186219 56897
rect 186247 56869 186281 56897
rect 186309 56869 201579 56897
rect 201607 56869 201641 56897
rect 201669 56869 216939 56897
rect 216967 56869 217001 56897
rect 217029 56869 232299 56897
rect 232327 56869 232361 56897
rect 232389 56869 247659 56897
rect 247687 56869 247721 56897
rect 247749 56869 254577 56897
rect 254605 56869 254639 56897
rect 254667 56869 254701 56897
rect 254729 56869 254763 56897
rect 254791 56869 263577 56897
rect 263605 56869 263639 56897
rect 263667 56869 263701 56897
rect 263729 56869 263763 56897
rect 263791 56869 272577 56897
rect 272605 56869 272639 56897
rect 272667 56869 272701 56897
rect 272729 56869 272763 56897
rect 272791 56869 281577 56897
rect 281605 56869 281639 56897
rect 281667 56869 281701 56897
rect 281729 56869 281763 56897
rect 281791 56869 290577 56897
rect 290605 56869 290639 56897
rect 290667 56869 290701 56897
rect 290729 56869 290763 56897
rect 290791 56869 299256 56897
rect 299284 56869 299318 56897
rect 299346 56869 299380 56897
rect 299408 56869 299442 56897
rect 299470 56869 299998 56897
rect -6 56835 299998 56869
rect -6 56807 522 56835
rect 550 56807 584 56835
rect 612 56807 646 56835
rect 674 56807 708 56835
rect 736 56807 2577 56835
rect 2605 56807 2639 56835
rect 2667 56807 2701 56835
rect 2729 56807 2763 56835
rect 2791 56807 11577 56835
rect 11605 56807 11639 56835
rect 11667 56807 11701 56835
rect 11729 56807 11763 56835
rect 11791 56807 17259 56835
rect 17287 56807 17321 56835
rect 17349 56807 20577 56835
rect 20605 56807 20639 56835
rect 20667 56807 20701 56835
rect 20729 56807 20763 56835
rect 20791 56807 29577 56835
rect 29605 56807 29639 56835
rect 29667 56807 29701 56835
rect 29729 56807 29763 56835
rect 29791 56807 32619 56835
rect 32647 56807 32681 56835
rect 32709 56807 47979 56835
rect 48007 56807 48041 56835
rect 48069 56807 63339 56835
rect 63367 56807 63401 56835
rect 63429 56807 78699 56835
rect 78727 56807 78761 56835
rect 78789 56807 94059 56835
rect 94087 56807 94121 56835
rect 94149 56807 109419 56835
rect 109447 56807 109481 56835
rect 109509 56807 124779 56835
rect 124807 56807 124841 56835
rect 124869 56807 140139 56835
rect 140167 56807 140201 56835
rect 140229 56807 155499 56835
rect 155527 56807 155561 56835
rect 155589 56807 170859 56835
rect 170887 56807 170921 56835
rect 170949 56807 186219 56835
rect 186247 56807 186281 56835
rect 186309 56807 201579 56835
rect 201607 56807 201641 56835
rect 201669 56807 216939 56835
rect 216967 56807 217001 56835
rect 217029 56807 232299 56835
rect 232327 56807 232361 56835
rect 232389 56807 247659 56835
rect 247687 56807 247721 56835
rect 247749 56807 254577 56835
rect 254605 56807 254639 56835
rect 254667 56807 254701 56835
rect 254729 56807 254763 56835
rect 254791 56807 263577 56835
rect 263605 56807 263639 56835
rect 263667 56807 263701 56835
rect 263729 56807 263763 56835
rect 263791 56807 272577 56835
rect 272605 56807 272639 56835
rect 272667 56807 272701 56835
rect 272729 56807 272763 56835
rect 272791 56807 281577 56835
rect 281605 56807 281639 56835
rect 281667 56807 281701 56835
rect 281729 56807 281763 56835
rect 281791 56807 290577 56835
rect 290605 56807 290639 56835
rect 290667 56807 290701 56835
rect 290729 56807 290763 56835
rect 290791 56807 299256 56835
rect 299284 56807 299318 56835
rect 299346 56807 299380 56835
rect 299408 56807 299442 56835
rect 299470 56807 299998 56835
rect -6 56773 299998 56807
rect -6 56745 522 56773
rect 550 56745 584 56773
rect 612 56745 646 56773
rect 674 56745 708 56773
rect 736 56745 2577 56773
rect 2605 56745 2639 56773
rect 2667 56745 2701 56773
rect 2729 56745 2763 56773
rect 2791 56745 11577 56773
rect 11605 56745 11639 56773
rect 11667 56745 11701 56773
rect 11729 56745 11763 56773
rect 11791 56745 17259 56773
rect 17287 56745 17321 56773
rect 17349 56745 20577 56773
rect 20605 56745 20639 56773
rect 20667 56745 20701 56773
rect 20729 56745 20763 56773
rect 20791 56745 29577 56773
rect 29605 56745 29639 56773
rect 29667 56745 29701 56773
rect 29729 56745 29763 56773
rect 29791 56745 32619 56773
rect 32647 56745 32681 56773
rect 32709 56745 47979 56773
rect 48007 56745 48041 56773
rect 48069 56745 63339 56773
rect 63367 56745 63401 56773
rect 63429 56745 78699 56773
rect 78727 56745 78761 56773
rect 78789 56745 94059 56773
rect 94087 56745 94121 56773
rect 94149 56745 109419 56773
rect 109447 56745 109481 56773
rect 109509 56745 124779 56773
rect 124807 56745 124841 56773
rect 124869 56745 140139 56773
rect 140167 56745 140201 56773
rect 140229 56745 155499 56773
rect 155527 56745 155561 56773
rect 155589 56745 170859 56773
rect 170887 56745 170921 56773
rect 170949 56745 186219 56773
rect 186247 56745 186281 56773
rect 186309 56745 201579 56773
rect 201607 56745 201641 56773
rect 201669 56745 216939 56773
rect 216967 56745 217001 56773
rect 217029 56745 232299 56773
rect 232327 56745 232361 56773
rect 232389 56745 247659 56773
rect 247687 56745 247721 56773
rect 247749 56745 254577 56773
rect 254605 56745 254639 56773
rect 254667 56745 254701 56773
rect 254729 56745 254763 56773
rect 254791 56745 263577 56773
rect 263605 56745 263639 56773
rect 263667 56745 263701 56773
rect 263729 56745 263763 56773
rect 263791 56745 272577 56773
rect 272605 56745 272639 56773
rect 272667 56745 272701 56773
rect 272729 56745 272763 56773
rect 272791 56745 281577 56773
rect 281605 56745 281639 56773
rect 281667 56745 281701 56773
rect 281729 56745 281763 56773
rect 281791 56745 290577 56773
rect 290605 56745 290639 56773
rect 290667 56745 290701 56773
rect 290729 56745 290763 56773
rect 290791 56745 299256 56773
rect 299284 56745 299318 56773
rect 299346 56745 299380 56773
rect 299408 56745 299442 56773
rect 299470 56745 299998 56773
rect -6 56697 299998 56745
rect -6 50959 299998 51007
rect -6 50931 42 50959
rect 70 50931 104 50959
rect 132 50931 166 50959
rect 194 50931 228 50959
rect 256 50931 4437 50959
rect 4465 50931 4499 50959
rect 4527 50931 4561 50959
rect 4589 50931 4623 50959
rect 4651 50931 13437 50959
rect 13465 50931 13499 50959
rect 13527 50931 13561 50959
rect 13589 50931 13623 50959
rect 13651 50931 22437 50959
rect 22465 50931 22499 50959
rect 22527 50931 22561 50959
rect 22589 50931 22623 50959
rect 22651 50931 24939 50959
rect 24967 50931 25001 50959
rect 25029 50931 31437 50959
rect 31465 50931 31499 50959
rect 31527 50931 31561 50959
rect 31589 50931 31623 50959
rect 31651 50931 40299 50959
rect 40327 50931 40361 50959
rect 40389 50931 55659 50959
rect 55687 50931 55721 50959
rect 55749 50931 71019 50959
rect 71047 50931 71081 50959
rect 71109 50931 86379 50959
rect 86407 50931 86441 50959
rect 86469 50931 101739 50959
rect 101767 50931 101801 50959
rect 101829 50931 117099 50959
rect 117127 50931 117161 50959
rect 117189 50931 132459 50959
rect 132487 50931 132521 50959
rect 132549 50931 147819 50959
rect 147847 50931 147881 50959
rect 147909 50931 163179 50959
rect 163207 50931 163241 50959
rect 163269 50931 178539 50959
rect 178567 50931 178601 50959
rect 178629 50931 193899 50959
rect 193927 50931 193961 50959
rect 193989 50931 209259 50959
rect 209287 50931 209321 50959
rect 209349 50931 224619 50959
rect 224647 50931 224681 50959
rect 224709 50931 239979 50959
rect 240007 50931 240041 50959
rect 240069 50931 256437 50959
rect 256465 50931 256499 50959
rect 256527 50931 256561 50959
rect 256589 50931 256623 50959
rect 256651 50931 265437 50959
rect 265465 50931 265499 50959
rect 265527 50931 265561 50959
rect 265589 50931 265623 50959
rect 265651 50931 274437 50959
rect 274465 50931 274499 50959
rect 274527 50931 274561 50959
rect 274589 50931 274623 50959
rect 274651 50931 283437 50959
rect 283465 50931 283499 50959
rect 283527 50931 283561 50959
rect 283589 50931 283623 50959
rect 283651 50931 292437 50959
rect 292465 50931 292499 50959
rect 292527 50931 292561 50959
rect 292589 50931 292623 50959
rect 292651 50931 299736 50959
rect 299764 50931 299798 50959
rect 299826 50931 299860 50959
rect 299888 50931 299922 50959
rect 299950 50931 299998 50959
rect -6 50897 299998 50931
rect -6 50869 42 50897
rect 70 50869 104 50897
rect 132 50869 166 50897
rect 194 50869 228 50897
rect 256 50869 4437 50897
rect 4465 50869 4499 50897
rect 4527 50869 4561 50897
rect 4589 50869 4623 50897
rect 4651 50869 13437 50897
rect 13465 50869 13499 50897
rect 13527 50869 13561 50897
rect 13589 50869 13623 50897
rect 13651 50869 22437 50897
rect 22465 50869 22499 50897
rect 22527 50869 22561 50897
rect 22589 50869 22623 50897
rect 22651 50869 24939 50897
rect 24967 50869 25001 50897
rect 25029 50869 31437 50897
rect 31465 50869 31499 50897
rect 31527 50869 31561 50897
rect 31589 50869 31623 50897
rect 31651 50869 40299 50897
rect 40327 50869 40361 50897
rect 40389 50869 55659 50897
rect 55687 50869 55721 50897
rect 55749 50869 71019 50897
rect 71047 50869 71081 50897
rect 71109 50869 86379 50897
rect 86407 50869 86441 50897
rect 86469 50869 101739 50897
rect 101767 50869 101801 50897
rect 101829 50869 117099 50897
rect 117127 50869 117161 50897
rect 117189 50869 132459 50897
rect 132487 50869 132521 50897
rect 132549 50869 147819 50897
rect 147847 50869 147881 50897
rect 147909 50869 163179 50897
rect 163207 50869 163241 50897
rect 163269 50869 178539 50897
rect 178567 50869 178601 50897
rect 178629 50869 193899 50897
rect 193927 50869 193961 50897
rect 193989 50869 209259 50897
rect 209287 50869 209321 50897
rect 209349 50869 224619 50897
rect 224647 50869 224681 50897
rect 224709 50869 239979 50897
rect 240007 50869 240041 50897
rect 240069 50869 256437 50897
rect 256465 50869 256499 50897
rect 256527 50869 256561 50897
rect 256589 50869 256623 50897
rect 256651 50869 265437 50897
rect 265465 50869 265499 50897
rect 265527 50869 265561 50897
rect 265589 50869 265623 50897
rect 265651 50869 274437 50897
rect 274465 50869 274499 50897
rect 274527 50869 274561 50897
rect 274589 50869 274623 50897
rect 274651 50869 283437 50897
rect 283465 50869 283499 50897
rect 283527 50869 283561 50897
rect 283589 50869 283623 50897
rect 283651 50869 292437 50897
rect 292465 50869 292499 50897
rect 292527 50869 292561 50897
rect 292589 50869 292623 50897
rect 292651 50869 299736 50897
rect 299764 50869 299798 50897
rect 299826 50869 299860 50897
rect 299888 50869 299922 50897
rect 299950 50869 299998 50897
rect -6 50835 299998 50869
rect -6 50807 42 50835
rect 70 50807 104 50835
rect 132 50807 166 50835
rect 194 50807 228 50835
rect 256 50807 4437 50835
rect 4465 50807 4499 50835
rect 4527 50807 4561 50835
rect 4589 50807 4623 50835
rect 4651 50807 13437 50835
rect 13465 50807 13499 50835
rect 13527 50807 13561 50835
rect 13589 50807 13623 50835
rect 13651 50807 22437 50835
rect 22465 50807 22499 50835
rect 22527 50807 22561 50835
rect 22589 50807 22623 50835
rect 22651 50807 24939 50835
rect 24967 50807 25001 50835
rect 25029 50807 31437 50835
rect 31465 50807 31499 50835
rect 31527 50807 31561 50835
rect 31589 50807 31623 50835
rect 31651 50807 40299 50835
rect 40327 50807 40361 50835
rect 40389 50807 55659 50835
rect 55687 50807 55721 50835
rect 55749 50807 71019 50835
rect 71047 50807 71081 50835
rect 71109 50807 86379 50835
rect 86407 50807 86441 50835
rect 86469 50807 101739 50835
rect 101767 50807 101801 50835
rect 101829 50807 117099 50835
rect 117127 50807 117161 50835
rect 117189 50807 132459 50835
rect 132487 50807 132521 50835
rect 132549 50807 147819 50835
rect 147847 50807 147881 50835
rect 147909 50807 163179 50835
rect 163207 50807 163241 50835
rect 163269 50807 178539 50835
rect 178567 50807 178601 50835
rect 178629 50807 193899 50835
rect 193927 50807 193961 50835
rect 193989 50807 209259 50835
rect 209287 50807 209321 50835
rect 209349 50807 224619 50835
rect 224647 50807 224681 50835
rect 224709 50807 239979 50835
rect 240007 50807 240041 50835
rect 240069 50807 256437 50835
rect 256465 50807 256499 50835
rect 256527 50807 256561 50835
rect 256589 50807 256623 50835
rect 256651 50807 265437 50835
rect 265465 50807 265499 50835
rect 265527 50807 265561 50835
rect 265589 50807 265623 50835
rect 265651 50807 274437 50835
rect 274465 50807 274499 50835
rect 274527 50807 274561 50835
rect 274589 50807 274623 50835
rect 274651 50807 283437 50835
rect 283465 50807 283499 50835
rect 283527 50807 283561 50835
rect 283589 50807 283623 50835
rect 283651 50807 292437 50835
rect 292465 50807 292499 50835
rect 292527 50807 292561 50835
rect 292589 50807 292623 50835
rect 292651 50807 299736 50835
rect 299764 50807 299798 50835
rect 299826 50807 299860 50835
rect 299888 50807 299922 50835
rect 299950 50807 299998 50835
rect -6 50773 299998 50807
rect -6 50745 42 50773
rect 70 50745 104 50773
rect 132 50745 166 50773
rect 194 50745 228 50773
rect 256 50745 4437 50773
rect 4465 50745 4499 50773
rect 4527 50745 4561 50773
rect 4589 50745 4623 50773
rect 4651 50745 13437 50773
rect 13465 50745 13499 50773
rect 13527 50745 13561 50773
rect 13589 50745 13623 50773
rect 13651 50745 22437 50773
rect 22465 50745 22499 50773
rect 22527 50745 22561 50773
rect 22589 50745 22623 50773
rect 22651 50745 24939 50773
rect 24967 50745 25001 50773
rect 25029 50745 31437 50773
rect 31465 50745 31499 50773
rect 31527 50745 31561 50773
rect 31589 50745 31623 50773
rect 31651 50745 40299 50773
rect 40327 50745 40361 50773
rect 40389 50745 55659 50773
rect 55687 50745 55721 50773
rect 55749 50745 71019 50773
rect 71047 50745 71081 50773
rect 71109 50745 86379 50773
rect 86407 50745 86441 50773
rect 86469 50745 101739 50773
rect 101767 50745 101801 50773
rect 101829 50745 117099 50773
rect 117127 50745 117161 50773
rect 117189 50745 132459 50773
rect 132487 50745 132521 50773
rect 132549 50745 147819 50773
rect 147847 50745 147881 50773
rect 147909 50745 163179 50773
rect 163207 50745 163241 50773
rect 163269 50745 178539 50773
rect 178567 50745 178601 50773
rect 178629 50745 193899 50773
rect 193927 50745 193961 50773
rect 193989 50745 209259 50773
rect 209287 50745 209321 50773
rect 209349 50745 224619 50773
rect 224647 50745 224681 50773
rect 224709 50745 239979 50773
rect 240007 50745 240041 50773
rect 240069 50745 256437 50773
rect 256465 50745 256499 50773
rect 256527 50745 256561 50773
rect 256589 50745 256623 50773
rect 256651 50745 265437 50773
rect 265465 50745 265499 50773
rect 265527 50745 265561 50773
rect 265589 50745 265623 50773
rect 265651 50745 274437 50773
rect 274465 50745 274499 50773
rect 274527 50745 274561 50773
rect 274589 50745 274623 50773
rect 274651 50745 283437 50773
rect 283465 50745 283499 50773
rect 283527 50745 283561 50773
rect 283589 50745 283623 50773
rect 283651 50745 292437 50773
rect 292465 50745 292499 50773
rect 292527 50745 292561 50773
rect 292589 50745 292623 50773
rect 292651 50745 299736 50773
rect 299764 50745 299798 50773
rect 299826 50745 299860 50773
rect 299888 50745 299922 50773
rect 299950 50745 299998 50773
rect -6 50697 299998 50745
rect -6 47959 299998 48007
rect -6 47931 522 47959
rect 550 47931 584 47959
rect 612 47931 646 47959
rect 674 47931 708 47959
rect 736 47931 2577 47959
rect 2605 47931 2639 47959
rect 2667 47931 2701 47959
rect 2729 47931 2763 47959
rect 2791 47931 11577 47959
rect 11605 47931 11639 47959
rect 11667 47931 11701 47959
rect 11729 47931 11763 47959
rect 11791 47931 17259 47959
rect 17287 47931 17321 47959
rect 17349 47931 20577 47959
rect 20605 47931 20639 47959
rect 20667 47931 20701 47959
rect 20729 47931 20763 47959
rect 20791 47931 29577 47959
rect 29605 47931 29639 47959
rect 29667 47931 29701 47959
rect 29729 47931 29763 47959
rect 29791 47931 32619 47959
rect 32647 47931 32681 47959
rect 32709 47931 47979 47959
rect 48007 47931 48041 47959
rect 48069 47931 63339 47959
rect 63367 47931 63401 47959
rect 63429 47931 78699 47959
rect 78727 47931 78761 47959
rect 78789 47931 94059 47959
rect 94087 47931 94121 47959
rect 94149 47931 109419 47959
rect 109447 47931 109481 47959
rect 109509 47931 124779 47959
rect 124807 47931 124841 47959
rect 124869 47931 140139 47959
rect 140167 47931 140201 47959
rect 140229 47931 155499 47959
rect 155527 47931 155561 47959
rect 155589 47931 170859 47959
rect 170887 47931 170921 47959
rect 170949 47931 186219 47959
rect 186247 47931 186281 47959
rect 186309 47931 201579 47959
rect 201607 47931 201641 47959
rect 201669 47931 216939 47959
rect 216967 47931 217001 47959
rect 217029 47931 232299 47959
rect 232327 47931 232361 47959
rect 232389 47931 247659 47959
rect 247687 47931 247721 47959
rect 247749 47931 254577 47959
rect 254605 47931 254639 47959
rect 254667 47931 254701 47959
rect 254729 47931 254763 47959
rect 254791 47931 263577 47959
rect 263605 47931 263639 47959
rect 263667 47931 263701 47959
rect 263729 47931 263763 47959
rect 263791 47931 272577 47959
rect 272605 47931 272639 47959
rect 272667 47931 272701 47959
rect 272729 47931 272763 47959
rect 272791 47931 281577 47959
rect 281605 47931 281639 47959
rect 281667 47931 281701 47959
rect 281729 47931 281763 47959
rect 281791 47931 290577 47959
rect 290605 47931 290639 47959
rect 290667 47931 290701 47959
rect 290729 47931 290763 47959
rect 290791 47931 299256 47959
rect 299284 47931 299318 47959
rect 299346 47931 299380 47959
rect 299408 47931 299442 47959
rect 299470 47931 299998 47959
rect -6 47897 299998 47931
rect -6 47869 522 47897
rect 550 47869 584 47897
rect 612 47869 646 47897
rect 674 47869 708 47897
rect 736 47869 2577 47897
rect 2605 47869 2639 47897
rect 2667 47869 2701 47897
rect 2729 47869 2763 47897
rect 2791 47869 11577 47897
rect 11605 47869 11639 47897
rect 11667 47869 11701 47897
rect 11729 47869 11763 47897
rect 11791 47869 17259 47897
rect 17287 47869 17321 47897
rect 17349 47869 20577 47897
rect 20605 47869 20639 47897
rect 20667 47869 20701 47897
rect 20729 47869 20763 47897
rect 20791 47869 29577 47897
rect 29605 47869 29639 47897
rect 29667 47869 29701 47897
rect 29729 47869 29763 47897
rect 29791 47869 32619 47897
rect 32647 47869 32681 47897
rect 32709 47869 47979 47897
rect 48007 47869 48041 47897
rect 48069 47869 63339 47897
rect 63367 47869 63401 47897
rect 63429 47869 78699 47897
rect 78727 47869 78761 47897
rect 78789 47869 94059 47897
rect 94087 47869 94121 47897
rect 94149 47869 109419 47897
rect 109447 47869 109481 47897
rect 109509 47869 124779 47897
rect 124807 47869 124841 47897
rect 124869 47869 140139 47897
rect 140167 47869 140201 47897
rect 140229 47869 155499 47897
rect 155527 47869 155561 47897
rect 155589 47869 170859 47897
rect 170887 47869 170921 47897
rect 170949 47869 186219 47897
rect 186247 47869 186281 47897
rect 186309 47869 201579 47897
rect 201607 47869 201641 47897
rect 201669 47869 216939 47897
rect 216967 47869 217001 47897
rect 217029 47869 232299 47897
rect 232327 47869 232361 47897
rect 232389 47869 247659 47897
rect 247687 47869 247721 47897
rect 247749 47869 254577 47897
rect 254605 47869 254639 47897
rect 254667 47869 254701 47897
rect 254729 47869 254763 47897
rect 254791 47869 263577 47897
rect 263605 47869 263639 47897
rect 263667 47869 263701 47897
rect 263729 47869 263763 47897
rect 263791 47869 272577 47897
rect 272605 47869 272639 47897
rect 272667 47869 272701 47897
rect 272729 47869 272763 47897
rect 272791 47869 281577 47897
rect 281605 47869 281639 47897
rect 281667 47869 281701 47897
rect 281729 47869 281763 47897
rect 281791 47869 290577 47897
rect 290605 47869 290639 47897
rect 290667 47869 290701 47897
rect 290729 47869 290763 47897
rect 290791 47869 299256 47897
rect 299284 47869 299318 47897
rect 299346 47869 299380 47897
rect 299408 47869 299442 47897
rect 299470 47869 299998 47897
rect -6 47835 299998 47869
rect -6 47807 522 47835
rect 550 47807 584 47835
rect 612 47807 646 47835
rect 674 47807 708 47835
rect 736 47807 2577 47835
rect 2605 47807 2639 47835
rect 2667 47807 2701 47835
rect 2729 47807 2763 47835
rect 2791 47807 11577 47835
rect 11605 47807 11639 47835
rect 11667 47807 11701 47835
rect 11729 47807 11763 47835
rect 11791 47807 17259 47835
rect 17287 47807 17321 47835
rect 17349 47807 20577 47835
rect 20605 47807 20639 47835
rect 20667 47807 20701 47835
rect 20729 47807 20763 47835
rect 20791 47807 29577 47835
rect 29605 47807 29639 47835
rect 29667 47807 29701 47835
rect 29729 47807 29763 47835
rect 29791 47807 32619 47835
rect 32647 47807 32681 47835
rect 32709 47807 47979 47835
rect 48007 47807 48041 47835
rect 48069 47807 63339 47835
rect 63367 47807 63401 47835
rect 63429 47807 78699 47835
rect 78727 47807 78761 47835
rect 78789 47807 94059 47835
rect 94087 47807 94121 47835
rect 94149 47807 109419 47835
rect 109447 47807 109481 47835
rect 109509 47807 124779 47835
rect 124807 47807 124841 47835
rect 124869 47807 140139 47835
rect 140167 47807 140201 47835
rect 140229 47807 155499 47835
rect 155527 47807 155561 47835
rect 155589 47807 170859 47835
rect 170887 47807 170921 47835
rect 170949 47807 186219 47835
rect 186247 47807 186281 47835
rect 186309 47807 201579 47835
rect 201607 47807 201641 47835
rect 201669 47807 216939 47835
rect 216967 47807 217001 47835
rect 217029 47807 232299 47835
rect 232327 47807 232361 47835
rect 232389 47807 247659 47835
rect 247687 47807 247721 47835
rect 247749 47807 254577 47835
rect 254605 47807 254639 47835
rect 254667 47807 254701 47835
rect 254729 47807 254763 47835
rect 254791 47807 263577 47835
rect 263605 47807 263639 47835
rect 263667 47807 263701 47835
rect 263729 47807 263763 47835
rect 263791 47807 272577 47835
rect 272605 47807 272639 47835
rect 272667 47807 272701 47835
rect 272729 47807 272763 47835
rect 272791 47807 281577 47835
rect 281605 47807 281639 47835
rect 281667 47807 281701 47835
rect 281729 47807 281763 47835
rect 281791 47807 290577 47835
rect 290605 47807 290639 47835
rect 290667 47807 290701 47835
rect 290729 47807 290763 47835
rect 290791 47807 299256 47835
rect 299284 47807 299318 47835
rect 299346 47807 299380 47835
rect 299408 47807 299442 47835
rect 299470 47807 299998 47835
rect -6 47773 299998 47807
rect -6 47745 522 47773
rect 550 47745 584 47773
rect 612 47745 646 47773
rect 674 47745 708 47773
rect 736 47745 2577 47773
rect 2605 47745 2639 47773
rect 2667 47745 2701 47773
rect 2729 47745 2763 47773
rect 2791 47745 11577 47773
rect 11605 47745 11639 47773
rect 11667 47745 11701 47773
rect 11729 47745 11763 47773
rect 11791 47745 17259 47773
rect 17287 47745 17321 47773
rect 17349 47745 20577 47773
rect 20605 47745 20639 47773
rect 20667 47745 20701 47773
rect 20729 47745 20763 47773
rect 20791 47745 29577 47773
rect 29605 47745 29639 47773
rect 29667 47745 29701 47773
rect 29729 47745 29763 47773
rect 29791 47745 32619 47773
rect 32647 47745 32681 47773
rect 32709 47745 47979 47773
rect 48007 47745 48041 47773
rect 48069 47745 63339 47773
rect 63367 47745 63401 47773
rect 63429 47745 78699 47773
rect 78727 47745 78761 47773
rect 78789 47745 94059 47773
rect 94087 47745 94121 47773
rect 94149 47745 109419 47773
rect 109447 47745 109481 47773
rect 109509 47745 124779 47773
rect 124807 47745 124841 47773
rect 124869 47745 140139 47773
rect 140167 47745 140201 47773
rect 140229 47745 155499 47773
rect 155527 47745 155561 47773
rect 155589 47745 170859 47773
rect 170887 47745 170921 47773
rect 170949 47745 186219 47773
rect 186247 47745 186281 47773
rect 186309 47745 201579 47773
rect 201607 47745 201641 47773
rect 201669 47745 216939 47773
rect 216967 47745 217001 47773
rect 217029 47745 232299 47773
rect 232327 47745 232361 47773
rect 232389 47745 247659 47773
rect 247687 47745 247721 47773
rect 247749 47745 254577 47773
rect 254605 47745 254639 47773
rect 254667 47745 254701 47773
rect 254729 47745 254763 47773
rect 254791 47745 263577 47773
rect 263605 47745 263639 47773
rect 263667 47745 263701 47773
rect 263729 47745 263763 47773
rect 263791 47745 272577 47773
rect 272605 47745 272639 47773
rect 272667 47745 272701 47773
rect 272729 47745 272763 47773
rect 272791 47745 281577 47773
rect 281605 47745 281639 47773
rect 281667 47745 281701 47773
rect 281729 47745 281763 47773
rect 281791 47745 290577 47773
rect 290605 47745 290639 47773
rect 290667 47745 290701 47773
rect 290729 47745 290763 47773
rect 290791 47745 299256 47773
rect 299284 47745 299318 47773
rect 299346 47745 299380 47773
rect 299408 47745 299442 47773
rect 299470 47745 299998 47773
rect -6 47697 299998 47745
rect -6 41959 299998 42007
rect -6 41931 42 41959
rect 70 41931 104 41959
rect 132 41931 166 41959
rect 194 41931 228 41959
rect 256 41931 4437 41959
rect 4465 41931 4499 41959
rect 4527 41931 4561 41959
rect 4589 41931 4623 41959
rect 4651 41931 13437 41959
rect 13465 41931 13499 41959
rect 13527 41931 13561 41959
rect 13589 41931 13623 41959
rect 13651 41931 22437 41959
rect 22465 41931 22499 41959
rect 22527 41931 22561 41959
rect 22589 41931 22623 41959
rect 22651 41931 24939 41959
rect 24967 41931 25001 41959
rect 25029 41931 31437 41959
rect 31465 41931 31499 41959
rect 31527 41931 31561 41959
rect 31589 41931 31623 41959
rect 31651 41931 40299 41959
rect 40327 41931 40361 41959
rect 40389 41931 55659 41959
rect 55687 41931 55721 41959
rect 55749 41931 71019 41959
rect 71047 41931 71081 41959
rect 71109 41931 86379 41959
rect 86407 41931 86441 41959
rect 86469 41931 101739 41959
rect 101767 41931 101801 41959
rect 101829 41931 117099 41959
rect 117127 41931 117161 41959
rect 117189 41931 132459 41959
rect 132487 41931 132521 41959
rect 132549 41931 147819 41959
rect 147847 41931 147881 41959
rect 147909 41931 163179 41959
rect 163207 41931 163241 41959
rect 163269 41931 178539 41959
rect 178567 41931 178601 41959
rect 178629 41931 193899 41959
rect 193927 41931 193961 41959
rect 193989 41931 209259 41959
rect 209287 41931 209321 41959
rect 209349 41931 224619 41959
rect 224647 41931 224681 41959
rect 224709 41931 239979 41959
rect 240007 41931 240041 41959
rect 240069 41931 256437 41959
rect 256465 41931 256499 41959
rect 256527 41931 256561 41959
rect 256589 41931 256623 41959
rect 256651 41931 265437 41959
rect 265465 41931 265499 41959
rect 265527 41931 265561 41959
rect 265589 41931 265623 41959
rect 265651 41931 274437 41959
rect 274465 41931 274499 41959
rect 274527 41931 274561 41959
rect 274589 41931 274623 41959
rect 274651 41931 283437 41959
rect 283465 41931 283499 41959
rect 283527 41931 283561 41959
rect 283589 41931 283623 41959
rect 283651 41931 292437 41959
rect 292465 41931 292499 41959
rect 292527 41931 292561 41959
rect 292589 41931 292623 41959
rect 292651 41931 299736 41959
rect 299764 41931 299798 41959
rect 299826 41931 299860 41959
rect 299888 41931 299922 41959
rect 299950 41931 299998 41959
rect -6 41897 299998 41931
rect -6 41869 42 41897
rect 70 41869 104 41897
rect 132 41869 166 41897
rect 194 41869 228 41897
rect 256 41869 4437 41897
rect 4465 41869 4499 41897
rect 4527 41869 4561 41897
rect 4589 41869 4623 41897
rect 4651 41869 13437 41897
rect 13465 41869 13499 41897
rect 13527 41869 13561 41897
rect 13589 41869 13623 41897
rect 13651 41869 22437 41897
rect 22465 41869 22499 41897
rect 22527 41869 22561 41897
rect 22589 41869 22623 41897
rect 22651 41869 24939 41897
rect 24967 41869 25001 41897
rect 25029 41869 31437 41897
rect 31465 41869 31499 41897
rect 31527 41869 31561 41897
rect 31589 41869 31623 41897
rect 31651 41869 40299 41897
rect 40327 41869 40361 41897
rect 40389 41869 55659 41897
rect 55687 41869 55721 41897
rect 55749 41869 71019 41897
rect 71047 41869 71081 41897
rect 71109 41869 86379 41897
rect 86407 41869 86441 41897
rect 86469 41869 101739 41897
rect 101767 41869 101801 41897
rect 101829 41869 117099 41897
rect 117127 41869 117161 41897
rect 117189 41869 132459 41897
rect 132487 41869 132521 41897
rect 132549 41869 147819 41897
rect 147847 41869 147881 41897
rect 147909 41869 163179 41897
rect 163207 41869 163241 41897
rect 163269 41869 178539 41897
rect 178567 41869 178601 41897
rect 178629 41869 193899 41897
rect 193927 41869 193961 41897
rect 193989 41869 209259 41897
rect 209287 41869 209321 41897
rect 209349 41869 224619 41897
rect 224647 41869 224681 41897
rect 224709 41869 239979 41897
rect 240007 41869 240041 41897
rect 240069 41869 256437 41897
rect 256465 41869 256499 41897
rect 256527 41869 256561 41897
rect 256589 41869 256623 41897
rect 256651 41869 265437 41897
rect 265465 41869 265499 41897
rect 265527 41869 265561 41897
rect 265589 41869 265623 41897
rect 265651 41869 274437 41897
rect 274465 41869 274499 41897
rect 274527 41869 274561 41897
rect 274589 41869 274623 41897
rect 274651 41869 283437 41897
rect 283465 41869 283499 41897
rect 283527 41869 283561 41897
rect 283589 41869 283623 41897
rect 283651 41869 292437 41897
rect 292465 41869 292499 41897
rect 292527 41869 292561 41897
rect 292589 41869 292623 41897
rect 292651 41869 299736 41897
rect 299764 41869 299798 41897
rect 299826 41869 299860 41897
rect 299888 41869 299922 41897
rect 299950 41869 299998 41897
rect -6 41835 299998 41869
rect -6 41807 42 41835
rect 70 41807 104 41835
rect 132 41807 166 41835
rect 194 41807 228 41835
rect 256 41807 4437 41835
rect 4465 41807 4499 41835
rect 4527 41807 4561 41835
rect 4589 41807 4623 41835
rect 4651 41807 13437 41835
rect 13465 41807 13499 41835
rect 13527 41807 13561 41835
rect 13589 41807 13623 41835
rect 13651 41807 22437 41835
rect 22465 41807 22499 41835
rect 22527 41807 22561 41835
rect 22589 41807 22623 41835
rect 22651 41807 24939 41835
rect 24967 41807 25001 41835
rect 25029 41807 31437 41835
rect 31465 41807 31499 41835
rect 31527 41807 31561 41835
rect 31589 41807 31623 41835
rect 31651 41807 40299 41835
rect 40327 41807 40361 41835
rect 40389 41807 55659 41835
rect 55687 41807 55721 41835
rect 55749 41807 71019 41835
rect 71047 41807 71081 41835
rect 71109 41807 86379 41835
rect 86407 41807 86441 41835
rect 86469 41807 101739 41835
rect 101767 41807 101801 41835
rect 101829 41807 117099 41835
rect 117127 41807 117161 41835
rect 117189 41807 132459 41835
rect 132487 41807 132521 41835
rect 132549 41807 147819 41835
rect 147847 41807 147881 41835
rect 147909 41807 163179 41835
rect 163207 41807 163241 41835
rect 163269 41807 178539 41835
rect 178567 41807 178601 41835
rect 178629 41807 193899 41835
rect 193927 41807 193961 41835
rect 193989 41807 209259 41835
rect 209287 41807 209321 41835
rect 209349 41807 224619 41835
rect 224647 41807 224681 41835
rect 224709 41807 239979 41835
rect 240007 41807 240041 41835
rect 240069 41807 256437 41835
rect 256465 41807 256499 41835
rect 256527 41807 256561 41835
rect 256589 41807 256623 41835
rect 256651 41807 265437 41835
rect 265465 41807 265499 41835
rect 265527 41807 265561 41835
rect 265589 41807 265623 41835
rect 265651 41807 274437 41835
rect 274465 41807 274499 41835
rect 274527 41807 274561 41835
rect 274589 41807 274623 41835
rect 274651 41807 283437 41835
rect 283465 41807 283499 41835
rect 283527 41807 283561 41835
rect 283589 41807 283623 41835
rect 283651 41807 292437 41835
rect 292465 41807 292499 41835
rect 292527 41807 292561 41835
rect 292589 41807 292623 41835
rect 292651 41807 299736 41835
rect 299764 41807 299798 41835
rect 299826 41807 299860 41835
rect 299888 41807 299922 41835
rect 299950 41807 299998 41835
rect -6 41773 299998 41807
rect -6 41745 42 41773
rect 70 41745 104 41773
rect 132 41745 166 41773
rect 194 41745 228 41773
rect 256 41745 4437 41773
rect 4465 41745 4499 41773
rect 4527 41745 4561 41773
rect 4589 41745 4623 41773
rect 4651 41745 13437 41773
rect 13465 41745 13499 41773
rect 13527 41745 13561 41773
rect 13589 41745 13623 41773
rect 13651 41745 22437 41773
rect 22465 41745 22499 41773
rect 22527 41745 22561 41773
rect 22589 41745 22623 41773
rect 22651 41745 24939 41773
rect 24967 41745 25001 41773
rect 25029 41745 31437 41773
rect 31465 41745 31499 41773
rect 31527 41745 31561 41773
rect 31589 41745 31623 41773
rect 31651 41745 40299 41773
rect 40327 41745 40361 41773
rect 40389 41745 55659 41773
rect 55687 41745 55721 41773
rect 55749 41745 71019 41773
rect 71047 41745 71081 41773
rect 71109 41745 86379 41773
rect 86407 41745 86441 41773
rect 86469 41745 101739 41773
rect 101767 41745 101801 41773
rect 101829 41745 117099 41773
rect 117127 41745 117161 41773
rect 117189 41745 132459 41773
rect 132487 41745 132521 41773
rect 132549 41745 147819 41773
rect 147847 41745 147881 41773
rect 147909 41745 163179 41773
rect 163207 41745 163241 41773
rect 163269 41745 178539 41773
rect 178567 41745 178601 41773
rect 178629 41745 193899 41773
rect 193927 41745 193961 41773
rect 193989 41745 209259 41773
rect 209287 41745 209321 41773
rect 209349 41745 224619 41773
rect 224647 41745 224681 41773
rect 224709 41745 239979 41773
rect 240007 41745 240041 41773
rect 240069 41745 256437 41773
rect 256465 41745 256499 41773
rect 256527 41745 256561 41773
rect 256589 41745 256623 41773
rect 256651 41745 265437 41773
rect 265465 41745 265499 41773
rect 265527 41745 265561 41773
rect 265589 41745 265623 41773
rect 265651 41745 274437 41773
rect 274465 41745 274499 41773
rect 274527 41745 274561 41773
rect 274589 41745 274623 41773
rect 274651 41745 283437 41773
rect 283465 41745 283499 41773
rect 283527 41745 283561 41773
rect 283589 41745 283623 41773
rect 283651 41745 292437 41773
rect 292465 41745 292499 41773
rect 292527 41745 292561 41773
rect 292589 41745 292623 41773
rect 292651 41745 299736 41773
rect 299764 41745 299798 41773
rect 299826 41745 299860 41773
rect 299888 41745 299922 41773
rect 299950 41745 299998 41773
rect -6 41697 299998 41745
rect -6 38959 299998 39007
rect -6 38931 522 38959
rect 550 38931 584 38959
rect 612 38931 646 38959
rect 674 38931 708 38959
rect 736 38931 2577 38959
rect 2605 38931 2639 38959
rect 2667 38931 2701 38959
rect 2729 38931 2763 38959
rect 2791 38931 11577 38959
rect 11605 38931 11639 38959
rect 11667 38931 11701 38959
rect 11729 38931 11763 38959
rect 11791 38931 17259 38959
rect 17287 38931 17321 38959
rect 17349 38931 20577 38959
rect 20605 38931 20639 38959
rect 20667 38931 20701 38959
rect 20729 38931 20763 38959
rect 20791 38931 29577 38959
rect 29605 38931 29639 38959
rect 29667 38931 29701 38959
rect 29729 38931 29763 38959
rect 29791 38931 32619 38959
rect 32647 38931 32681 38959
rect 32709 38931 47979 38959
rect 48007 38931 48041 38959
rect 48069 38931 63339 38959
rect 63367 38931 63401 38959
rect 63429 38931 78699 38959
rect 78727 38931 78761 38959
rect 78789 38931 94059 38959
rect 94087 38931 94121 38959
rect 94149 38931 109419 38959
rect 109447 38931 109481 38959
rect 109509 38931 124779 38959
rect 124807 38931 124841 38959
rect 124869 38931 140139 38959
rect 140167 38931 140201 38959
rect 140229 38931 155499 38959
rect 155527 38931 155561 38959
rect 155589 38931 170859 38959
rect 170887 38931 170921 38959
rect 170949 38931 186219 38959
rect 186247 38931 186281 38959
rect 186309 38931 201579 38959
rect 201607 38931 201641 38959
rect 201669 38931 216939 38959
rect 216967 38931 217001 38959
rect 217029 38931 232299 38959
rect 232327 38931 232361 38959
rect 232389 38931 247659 38959
rect 247687 38931 247721 38959
rect 247749 38931 254577 38959
rect 254605 38931 254639 38959
rect 254667 38931 254701 38959
rect 254729 38931 254763 38959
rect 254791 38931 263577 38959
rect 263605 38931 263639 38959
rect 263667 38931 263701 38959
rect 263729 38931 263763 38959
rect 263791 38931 272577 38959
rect 272605 38931 272639 38959
rect 272667 38931 272701 38959
rect 272729 38931 272763 38959
rect 272791 38931 281577 38959
rect 281605 38931 281639 38959
rect 281667 38931 281701 38959
rect 281729 38931 281763 38959
rect 281791 38931 290577 38959
rect 290605 38931 290639 38959
rect 290667 38931 290701 38959
rect 290729 38931 290763 38959
rect 290791 38931 299256 38959
rect 299284 38931 299318 38959
rect 299346 38931 299380 38959
rect 299408 38931 299442 38959
rect 299470 38931 299998 38959
rect -6 38897 299998 38931
rect -6 38869 522 38897
rect 550 38869 584 38897
rect 612 38869 646 38897
rect 674 38869 708 38897
rect 736 38869 2577 38897
rect 2605 38869 2639 38897
rect 2667 38869 2701 38897
rect 2729 38869 2763 38897
rect 2791 38869 11577 38897
rect 11605 38869 11639 38897
rect 11667 38869 11701 38897
rect 11729 38869 11763 38897
rect 11791 38869 17259 38897
rect 17287 38869 17321 38897
rect 17349 38869 20577 38897
rect 20605 38869 20639 38897
rect 20667 38869 20701 38897
rect 20729 38869 20763 38897
rect 20791 38869 29577 38897
rect 29605 38869 29639 38897
rect 29667 38869 29701 38897
rect 29729 38869 29763 38897
rect 29791 38869 32619 38897
rect 32647 38869 32681 38897
rect 32709 38869 47979 38897
rect 48007 38869 48041 38897
rect 48069 38869 63339 38897
rect 63367 38869 63401 38897
rect 63429 38869 78699 38897
rect 78727 38869 78761 38897
rect 78789 38869 94059 38897
rect 94087 38869 94121 38897
rect 94149 38869 109419 38897
rect 109447 38869 109481 38897
rect 109509 38869 124779 38897
rect 124807 38869 124841 38897
rect 124869 38869 140139 38897
rect 140167 38869 140201 38897
rect 140229 38869 155499 38897
rect 155527 38869 155561 38897
rect 155589 38869 170859 38897
rect 170887 38869 170921 38897
rect 170949 38869 186219 38897
rect 186247 38869 186281 38897
rect 186309 38869 201579 38897
rect 201607 38869 201641 38897
rect 201669 38869 216939 38897
rect 216967 38869 217001 38897
rect 217029 38869 232299 38897
rect 232327 38869 232361 38897
rect 232389 38869 247659 38897
rect 247687 38869 247721 38897
rect 247749 38869 254577 38897
rect 254605 38869 254639 38897
rect 254667 38869 254701 38897
rect 254729 38869 254763 38897
rect 254791 38869 263577 38897
rect 263605 38869 263639 38897
rect 263667 38869 263701 38897
rect 263729 38869 263763 38897
rect 263791 38869 272577 38897
rect 272605 38869 272639 38897
rect 272667 38869 272701 38897
rect 272729 38869 272763 38897
rect 272791 38869 281577 38897
rect 281605 38869 281639 38897
rect 281667 38869 281701 38897
rect 281729 38869 281763 38897
rect 281791 38869 290577 38897
rect 290605 38869 290639 38897
rect 290667 38869 290701 38897
rect 290729 38869 290763 38897
rect 290791 38869 299256 38897
rect 299284 38869 299318 38897
rect 299346 38869 299380 38897
rect 299408 38869 299442 38897
rect 299470 38869 299998 38897
rect -6 38835 299998 38869
rect -6 38807 522 38835
rect 550 38807 584 38835
rect 612 38807 646 38835
rect 674 38807 708 38835
rect 736 38807 2577 38835
rect 2605 38807 2639 38835
rect 2667 38807 2701 38835
rect 2729 38807 2763 38835
rect 2791 38807 11577 38835
rect 11605 38807 11639 38835
rect 11667 38807 11701 38835
rect 11729 38807 11763 38835
rect 11791 38807 17259 38835
rect 17287 38807 17321 38835
rect 17349 38807 20577 38835
rect 20605 38807 20639 38835
rect 20667 38807 20701 38835
rect 20729 38807 20763 38835
rect 20791 38807 29577 38835
rect 29605 38807 29639 38835
rect 29667 38807 29701 38835
rect 29729 38807 29763 38835
rect 29791 38807 32619 38835
rect 32647 38807 32681 38835
rect 32709 38807 47979 38835
rect 48007 38807 48041 38835
rect 48069 38807 63339 38835
rect 63367 38807 63401 38835
rect 63429 38807 78699 38835
rect 78727 38807 78761 38835
rect 78789 38807 94059 38835
rect 94087 38807 94121 38835
rect 94149 38807 109419 38835
rect 109447 38807 109481 38835
rect 109509 38807 124779 38835
rect 124807 38807 124841 38835
rect 124869 38807 140139 38835
rect 140167 38807 140201 38835
rect 140229 38807 155499 38835
rect 155527 38807 155561 38835
rect 155589 38807 170859 38835
rect 170887 38807 170921 38835
rect 170949 38807 186219 38835
rect 186247 38807 186281 38835
rect 186309 38807 201579 38835
rect 201607 38807 201641 38835
rect 201669 38807 216939 38835
rect 216967 38807 217001 38835
rect 217029 38807 232299 38835
rect 232327 38807 232361 38835
rect 232389 38807 247659 38835
rect 247687 38807 247721 38835
rect 247749 38807 254577 38835
rect 254605 38807 254639 38835
rect 254667 38807 254701 38835
rect 254729 38807 254763 38835
rect 254791 38807 263577 38835
rect 263605 38807 263639 38835
rect 263667 38807 263701 38835
rect 263729 38807 263763 38835
rect 263791 38807 272577 38835
rect 272605 38807 272639 38835
rect 272667 38807 272701 38835
rect 272729 38807 272763 38835
rect 272791 38807 281577 38835
rect 281605 38807 281639 38835
rect 281667 38807 281701 38835
rect 281729 38807 281763 38835
rect 281791 38807 290577 38835
rect 290605 38807 290639 38835
rect 290667 38807 290701 38835
rect 290729 38807 290763 38835
rect 290791 38807 299256 38835
rect 299284 38807 299318 38835
rect 299346 38807 299380 38835
rect 299408 38807 299442 38835
rect 299470 38807 299998 38835
rect -6 38773 299998 38807
rect -6 38745 522 38773
rect 550 38745 584 38773
rect 612 38745 646 38773
rect 674 38745 708 38773
rect 736 38745 2577 38773
rect 2605 38745 2639 38773
rect 2667 38745 2701 38773
rect 2729 38745 2763 38773
rect 2791 38745 11577 38773
rect 11605 38745 11639 38773
rect 11667 38745 11701 38773
rect 11729 38745 11763 38773
rect 11791 38745 17259 38773
rect 17287 38745 17321 38773
rect 17349 38745 20577 38773
rect 20605 38745 20639 38773
rect 20667 38745 20701 38773
rect 20729 38745 20763 38773
rect 20791 38745 29577 38773
rect 29605 38745 29639 38773
rect 29667 38745 29701 38773
rect 29729 38745 29763 38773
rect 29791 38745 32619 38773
rect 32647 38745 32681 38773
rect 32709 38745 47979 38773
rect 48007 38745 48041 38773
rect 48069 38745 63339 38773
rect 63367 38745 63401 38773
rect 63429 38745 78699 38773
rect 78727 38745 78761 38773
rect 78789 38745 94059 38773
rect 94087 38745 94121 38773
rect 94149 38745 109419 38773
rect 109447 38745 109481 38773
rect 109509 38745 124779 38773
rect 124807 38745 124841 38773
rect 124869 38745 140139 38773
rect 140167 38745 140201 38773
rect 140229 38745 155499 38773
rect 155527 38745 155561 38773
rect 155589 38745 170859 38773
rect 170887 38745 170921 38773
rect 170949 38745 186219 38773
rect 186247 38745 186281 38773
rect 186309 38745 201579 38773
rect 201607 38745 201641 38773
rect 201669 38745 216939 38773
rect 216967 38745 217001 38773
rect 217029 38745 232299 38773
rect 232327 38745 232361 38773
rect 232389 38745 247659 38773
rect 247687 38745 247721 38773
rect 247749 38745 254577 38773
rect 254605 38745 254639 38773
rect 254667 38745 254701 38773
rect 254729 38745 254763 38773
rect 254791 38745 263577 38773
rect 263605 38745 263639 38773
rect 263667 38745 263701 38773
rect 263729 38745 263763 38773
rect 263791 38745 272577 38773
rect 272605 38745 272639 38773
rect 272667 38745 272701 38773
rect 272729 38745 272763 38773
rect 272791 38745 281577 38773
rect 281605 38745 281639 38773
rect 281667 38745 281701 38773
rect 281729 38745 281763 38773
rect 281791 38745 290577 38773
rect 290605 38745 290639 38773
rect 290667 38745 290701 38773
rect 290729 38745 290763 38773
rect 290791 38745 299256 38773
rect 299284 38745 299318 38773
rect 299346 38745 299380 38773
rect 299408 38745 299442 38773
rect 299470 38745 299998 38773
rect -6 38697 299998 38745
rect -6 32959 299998 33007
rect -6 32931 42 32959
rect 70 32931 104 32959
rect 132 32931 166 32959
rect 194 32931 228 32959
rect 256 32931 4437 32959
rect 4465 32931 4499 32959
rect 4527 32931 4561 32959
rect 4589 32931 4623 32959
rect 4651 32931 13437 32959
rect 13465 32931 13499 32959
rect 13527 32931 13561 32959
rect 13589 32931 13623 32959
rect 13651 32931 22437 32959
rect 22465 32931 22499 32959
rect 22527 32931 22561 32959
rect 22589 32931 22623 32959
rect 22651 32931 24939 32959
rect 24967 32931 25001 32959
rect 25029 32931 31437 32959
rect 31465 32931 31499 32959
rect 31527 32931 31561 32959
rect 31589 32931 31623 32959
rect 31651 32931 40299 32959
rect 40327 32931 40361 32959
rect 40389 32931 55659 32959
rect 55687 32931 55721 32959
rect 55749 32931 71019 32959
rect 71047 32931 71081 32959
rect 71109 32931 86379 32959
rect 86407 32931 86441 32959
rect 86469 32931 101739 32959
rect 101767 32931 101801 32959
rect 101829 32931 117099 32959
rect 117127 32931 117161 32959
rect 117189 32931 132459 32959
rect 132487 32931 132521 32959
rect 132549 32931 147819 32959
rect 147847 32931 147881 32959
rect 147909 32931 163179 32959
rect 163207 32931 163241 32959
rect 163269 32931 178539 32959
rect 178567 32931 178601 32959
rect 178629 32931 193899 32959
rect 193927 32931 193961 32959
rect 193989 32931 209259 32959
rect 209287 32931 209321 32959
rect 209349 32931 224619 32959
rect 224647 32931 224681 32959
rect 224709 32931 239979 32959
rect 240007 32931 240041 32959
rect 240069 32931 256437 32959
rect 256465 32931 256499 32959
rect 256527 32931 256561 32959
rect 256589 32931 256623 32959
rect 256651 32931 265437 32959
rect 265465 32931 265499 32959
rect 265527 32931 265561 32959
rect 265589 32931 265623 32959
rect 265651 32931 274437 32959
rect 274465 32931 274499 32959
rect 274527 32931 274561 32959
rect 274589 32931 274623 32959
rect 274651 32931 283437 32959
rect 283465 32931 283499 32959
rect 283527 32931 283561 32959
rect 283589 32931 283623 32959
rect 283651 32931 292437 32959
rect 292465 32931 292499 32959
rect 292527 32931 292561 32959
rect 292589 32931 292623 32959
rect 292651 32931 299736 32959
rect 299764 32931 299798 32959
rect 299826 32931 299860 32959
rect 299888 32931 299922 32959
rect 299950 32931 299998 32959
rect -6 32897 299998 32931
rect -6 32869 42 32897
rect 70 32869 104 32897
rect 132 32869 166 32897
rect 194 32869 228 32897
rect 256 32869 4437 32897
rect 4465 32869 4499 32897
rect 4527 32869 4561 32897
rect 4589 32869 4623 32897
rect 4651 32869 13437 32897
rect 13465 32869 13499 32897
rect 13527 32869 13561 32897
rect 13589 32869 13623 32897
rect 13651 32869 22437 32897
rect 22465 32869 22499 32897
rect 22527 32869 22561 32897
rect 22589 32869 22623 32897
rect 22651 32869 24939 32897
rect 24967 32869 25001 32897
rect 25029 32869 31437 32897
rect 31465 32869 31499 32897
rect 31527 32869 31561 32897
rect 31589 32869 31623 32897
rect 31651 32869 40299 32897
rect 40327 32869 40361 32897
rect 40389 32869 55659 32897
rect 55687 32869 55721 32897
rect 55749 32869 71019 32897
rect 71047 32869 71081 32897
rect 71109 32869 86379 32897
rect 86407 32869 86441 32897
rect 86469 32869 101739 32897
rect 101767 32869 101801 32897
rect 101829 32869 117099 32897
rect 117127 32869 117161 32897
rect 117189 32869 132459 32897
rect 132487 32869 132521 32897
rect 132549 32869 147819 32897
rect 147847 32869 147881 32897
rect 147909 32869 163179 32897
rect 163207 32869 163241 32897
rect 163269 32869 178539 32897
rect 178567 32869 178601 32897
rect 178629 32869 193899 32897
rect 193927 32869 193961 32897
rect 193989 32869 209259 32897
rect 209287 32869 209321 32897
rect 209349 32869 224619 32897
rect 224647 32869 224681 32897
rect 224709 32869 239979 32897
rect 240007 32869 240041 32897
rect 240069 32869 256437 32897
rect 256465 32869 256499 32897
rect 256527 32869 256561 32897
rect 256589 32869 256623 32897
rect 256651 32869 265437 32897
rect 265465 32869 265499 32897
rect 265527 32869 265561 32897
rect 265589 32869 265623 32897
rect 265651 32869 274437 32897
rect 274465 32869 274499 32897
rect 274527 32869 274561 32897
rect 274589 32869 274623 32897
rect 274651 32869 283437 32897
rect 283465 32869 283499 32897
rect 283527 32869 283561 32897
rect 283589 32869 283623 32897
rect 283651 32869 292437 32897
rect 292465 32869 292499 32897
rect 292527 32869 292561 32897
rect 292589 32869 292623 32897
rect 292651 32869 299736 32897
rect 299764 32869 299798 32897
rect 299826 32869 299860 32897
rect 299888 32869 299922 32897
rect 299950 32869 299998 32897
rect -6 32835 299998 32869
rect -6 32807 42 32835
rect 70 32807 104 32835
rect 132 32807 166 32835
rect 194 32807 228 32835
rect 256 32807 4437 32835
rect 4465 32807 4499 32835
rect 4527 32807 4561 32835
rect 4589 32807 4623 32835
rect 4651 32807 13437 32835
rect 13465 32807 13499 32835
rect 13527 32807 13561 32835
rect 13589 32807 13623 32835
rect 13651 32807 22437 32835
rect 22465 32807 22499 32835
rect 22527 32807 22561 32835
rect 22589 32807 22623 32835
rect 22651 32807 24939 32835
rect 24967 32807 25001 32835
rect 25029 32807 31437 32835
rect 31465 32807 31499 32835
rect 31527 32807 31561 32835
rect 31589 32807 31623 32835
rect 31651 32807 40299 32835
rect 40327 32807 40361 32835
rect 40389 32807 55659 32835
rect 55687 32807 55721 32835
rect 55749 32807 71019 32835
rect 71047 32807 71081 32835
rect 71109 32807 86379 32835
rect 86407 32807 86441 32835
rect 86469 32807 101739 32835
rect 101767 32807 101801 32835
rect 101829 32807 117099 32835
rect 117127 32807 117161 32835
rect 117189 32807 132459 32835
rect 132487 32807 132521 32835
rect 132549 32807 147819 32835
rect 147847 32807 147881 32835
rect 147909 32807 163179 32835
rect 163207 32807 163241 32835
rect 163269 32807 178539 32835
rect 178567 32807 178601 32835
rect 178629 32807 193899 32835
rect 193927 32807 193961 32835
rect 193989 32807 209259 32835
rect 209287 32807 209321 32835
rect 209349 32807 224619 32835
rect 224647 32807 224681 32835
rect 224709 32807 239979 32835
rect 240007 32807 240041 32835
rect 240069 32807 256437 32835
rect 256465 32807 256499 32835
rect 256527 32807 256561 32835
rect 256589 32807 256623 32835
rect 256651 32807 265437 32835
rect 265465 32807 265499 32835
rect 265527 32807 265561 32835
rect 265589 32807 265623 32835
rect 265651 32807 274437 32835
rect 274465 32807 274499 32835
rect 274527 32807 274561 32835
rect 274589 32807 274623 32835
rect 274651 32807 283437 32835
rect 283465 32807 283499 32835
rect 283527 32807 283561 32835
rect 283589 32807 283623 32835
rect 283651 32807 292437 32835
rect 292465 32807 292499 32835
rect 292527 32807 292561 32835
rect 292589 32807 292623 32835
rect 292651 32807 299736 32835
rect 299764 32807 299798 32835
rect 299826 32807 299860 32835
rect 299888 32807 299922 32835
rect 299950 32807 299998 32835
rect -6 32773 299998 32807
rect -6 32745 42 32773
rect 70 32745 104 32773
rect 132 32745 166 32773
rect 194 32745 228 32773
rect 256 32745 4437 32773
rect 4465 32745 4499 32773
rect 4527 32745 4561 32773
rect 4589 32745 4623 32773
rect 4651 32745 13437 32773
rect 13465 32745 13499 32773
rect 13527 32745 13561 32773
rect 13589 32745 13623 32773
rect 13651 32745 22437 32773
rect 22465 32745 22499 32773
rect 22527 32745 22561 32773
rect 22589 32745 22623 32773
rect 22651 32745 24939 32773
rect 24967 32745 25001 32773
rect 25029 32745 31437 32773
rect 31465 32745 31499 32773
rect 31527 32745 31561 32773
rect 31589 32745 31623 32773
rect 31651 32745 40299 32773
rect 40327 32745 40361 32773
rect 40389 32745 55659 32773
rect 55687 32745 55721 32773
rect 55749 32745 71019 32773
rect 71047 32745 71081 32773
rect 71109 32745 86379 32773
rect 86407 32745 86441 32773
rect 86469 32745 101739 32773
rect 101767 32745 101801 32773
rect 101829 32745 117099 32773
rect 117127 32745 117161 32773
rect 117189 32745 132459 32773
rect 132487 32745 132521 32773
rect 132549 32745 147819 32773
rect 147847 32745 147881 32773
rect 147909 32745 163179 32773
rect 163207 32745 163241 32773
rect 163269 32745 178539 32773
rect 178567 32745 178601 32773
rect 178629 32745 193899 32773
rect 193927 32745 193961 32773
rect 193989 32745 209259 32773
rect 209287 32745 209321 32773
rect 209349 32745 224619 32773
rect 224647 32745 224681 32773
rect 224709 32745 239979 32773
rect 240007 32745 240041 32773
rect 240069 32745 256437 32773
rect 256465 32745 256499 32773
rect 256527 32745 256561 32773
rect 256589 32745 256623 32773
rect 256651 32745 265437 32773
rect 265465 32745 265499 32773
rect 265527 32745 265561 32773
rect 265589 32745 265623 32773
rect 265651 32745 274437 32773
rect 274465 32745 274499 32773
rect 274527 32745 274561 32773
rect 274589 32745 274623 32773
rect 274651 32745 283437 32773
rect 283465 32745 283499 32773
rect 283527 32745 283561 32773
rect 283589 32745 283623 32773
rect 283651 32745 292437 32773
rect 292465 32745 292499 32773
rect 292527 32745 292561 32773
rect 292589 32745 292623 32773
rect 292651 32745 299736 32773
rect 299764 32745 299798 32773
rect 299826 32745 299860 32773
rect 299888 32745 299922 32773
rect 299950 32745 299998 32773
rect -6 32697 299998 32745
rect -6 29959 299998 30007
rect -6 29931 522 29959
rect 550 29931 584 29959
rect 612 29931 646 29959
rect 674 29931 708 29959
rect 736 29931 2577 29959
rect 2605 29931 2639 29959
rect 2667 29931 2701 29959
rect 2729 29931 2763 29959
rect 2791 29931 11577 29959
rect 11605 29931 11639 29959
rect 11667 29931 11701 29959
rect 11729 29931 11763 29959
rect 11791 29931 17259 29959
rect 17287 29931 17321 29959
rect 17349 29931 20577 29959
rect 20605 29931 20639 29959
rect 20667 29931 20701 29959
rect 20729 29931 20763 29959
rect 20791 29931 29577 29959
rect 29605 29931 29639 29959
rect 29667 29931 29701 29959
rect 29729 29931 29763 29959
rect 29791 29931 32619 29959
rect 32647 29931 32681 29959
rect 32709 29931 47979 29959
rect 48007 29931 48041 29959
rect 48069 29931 63339 29959
rect 63367 29931 63401 29959
rect 63429 29931 78699 29959
rect 78727 29931 78761 29959
rect 78789 29931 94059 29959
rect 94087 29931 94121 29959
rect 94149 29931 109419 29959
rect 109447 29931 109481 29959
rect 109509 29931 124779 29959
rect 124807 29931 124841 29959
rect 124869 29931 140139 29959
rect 140167 29931 140201 29959
rect 140229 29931 155499 29959
rect 155527 29931 155561 29959
rect 155589 29931 170859 29959
rect 170887 29931 170921 29959
rect 170949 29931 186219 29959
rect 186247 29931 186281 29959
rect 186309 29931 201579 29959
rect 201607 29931 201641 29959
rect 201669 29931 216939 29959
rect 216967 29931 217001 29959
rect 217029 29931 232299 29959
rect 232327 29931 232361 29959
rect 232389 29931 247659 29959
rect 247687 29931 247721 29959
rect 247749 29931 254577 29959
rect 254605 29931 254639 29959
rect 254667 29931 254701 29959
rect 254729 29931 254763 29959
rect 254791 29931 263577 29959
rect 263605 29931 263639 29959
rect 263667 29931 263701 29959
rect 263729 29931 263763 29959
rect 263791 29931 272577 29959
rect 272605 29931 272639 29959
rect 272667 29931 272701 29959
rect 272729 29931 272763 29959
rect 272791 29931 281577 29959
rect 281605 29931 281639 29959
rect 281667 29931 281701 29959
rect 281729 29931 281763 29959
rect 281791 29931 290577 29959
rect 290605 29931 290639 29959
rect 290667 29931 290701 29959
rect 290729 29931 290763 29959
rect 290791 29931 299256 29959
rect 299284 29931 299318 29959
rect 299346 29931 299380 29959
rect 299408 29931 299442 29959
rect 299470 29931 299998 29959
rect -6 29897 299998 29931
rect -6 29869 522 29897
rect 550 29869 584 29897
rect 612 29869 646 29897
rect 674 29869 708 29897
rect 736 29869 2577 29897
rect 2605 29869 2639 29897
rect 2667 29869 2701 29897
rect 2729 29869 2763 29897
rect 2791 29869 11577 29897
rect 11605 29869 11639 29897
rect 11667 29869 11701 29897
rect 11729 29869 11763 29897
rect 11791 29869 17259 29897
rect 17287 29869 17321 29897
rect 17349 29869 20577 29897
rect 20605 29869 20639 29897
rect 20667 29869 20701 29897
rect 20729 29869 20763 29897
rect 20791 29869 29577 29897
rect 29605 29869 29639 29897
rect 29667 29869 29701 29897
rect 29729 29869 29763 29897
rect 29791 29869 32619 29897
rect 32647 29869 32681 29897
rect 32709 29869 47979 29897
rect 48007 29869 48041 29897
rect 48069 29869 63339 29897
rect 63367 29869 63401 29897
rect 63429 29869 78699 29897
rect 78727 29869 78761 29897
rect 78789 29869 94059 29897
rect 94087 29869 94121 29897
rect 94149 29869 109419 29897
rect 109447 29869 109481 29897
rect 109509 29869 124779 29897
rect 124807 29869 124841 29897
rect 124869 29869 140139 29897
rect 140167 29869 140201 29897
rect 140229 29869 155499 29897
rect 155527 29869 155561 29897
rect 155589 29869 170859 29897
rect 170887 29869 170921 29897
rect 170949 29869 186219 29897
rect 186247 29869 186281 29897
rect 186309 29869 201579 29897
rect 201607 29869 201641 29897
rect 201669 29869 216939 29897
rect 216967 29869 217001 29897
rect 217029 29869 232299 29897
rect 232327 29869 232361 29897
rect 232389 29869 247659 29897
rect 247687 29869 247721 29897
rect 247749 29869 254577 29897
rect 254605 29869 254639 29897
rect 254667 29869 254701 29897
rect 254729 29869 254763 29897
rect 254791 29869 263577 29897
rect 263605 29869 263639 29897
rect 263667 29869 263701 29897
rect 263729 29869 263763 29897
rect 263791 29869 272577 29897
rect 272605 29869 272639 29897
rect 272667 29869 272701 29897
rect 272729 29869 272763 29897
rect 272791 29869 281577 29897
rect 281605 29869 281639 29897
rect 281667 29869 281701 29897
rect 281729 29869 281763 29897
rect 281791 29869 290577 29897
rect 290605 29869 290639 29897
rect 290667 29869 290701 29897
rect 290729 29869 290763 29897
rect 290791 29869 299256 29897
rect 299284 29869 299318 29897
rect 299346 29869 299380 29897
rect 299408 29869 299442 29897
rect 299470 29869 299998 29897
rect -6 29835 299998 29869
rect -6 29807 522 29835
rect 550 29807 584 29835
rect 612 29807 646 29835
rect 674 29807 708 29835
rect 736 29807 2577 29835
rect 2605 29807 2639 29835
rect 2667 29807 2701 29835
rect 2729 29807 2763 29835
rect 2791 29807 11577 29835
rect 11605 29807 11639 29835
rect 11667 29807 11701 29835
rect 11729 29807 11763 29835
rect 11791 29807 17259 29835
rect 17287 29807 17321 29835
rect 17349 29807 20577 29835
rect 20605 29807 20639 29835
rect 20667 29807 20701 29835
rect 20729 29807 20763 29835
rect 20791 29807 29577 29835
rect 29605 29807 29639 29835
rect 29667 29807 29701 29835
rect 29729 29807 29763 29835
rect 29791 29807 32619 29835
rect 32647 29807 32681 29835
rect 32709 29807 47979 29835
rect 48007 29807 48041 29835
rect 48069 29807 63339 29835
rect 63367 29807 63401 29835
rect 63429 29807 78699 29835
rect 78727 29807 78761 29835
rect 78789 29807 94059 29835
rect 94087 29807 94121 29835
rect 94149 29807 109419 29835
rect 109447 29807 109481 29835
rect 109509 29807 124779 29835
rect 124807 29807 124841 29835
rect 124869 29807 140139 29835
rect 140167 29807 140201 29835
rect 140229 29807 155499 29835
rect 155527 29807 155561 29835
rect 155589 29807 170859 29835
rect 170887 29807 170921 29835
rect 170949 29807 186219 29835
rect 186247 29807 186281 29835
rect 186309 29807 201579 29835
rect 201607 29807 201641 29835
rect 201669 29807 216939 29835
rect 216967 29807 217001 29835
rect 217029 29807 232299 29835
rect 232327 29807 232361 29835
rect 232389 29807 247659 29835
rect 247687 29807 247721 29835
rect 247749 29807 254577 29835
rect 254605 29807 254639 29835
rect 254667 29807 254701 29835
rect 254729 29807 254763 29835
rect 254791 29807 263577 29835
rect 263605 29807 263639 29835
rect 263667 29807 263701 29835
rect 263729 29807 263763 29835
rect 263791 29807 272577 29835
rect 272605 29807 272639 29835
rect 272667 29807 272701 29835
rect 272729 29807 272763 29835
rect 272791 29807 281577 29835
rect 281605 29807 281639 29835
rect 281667 29807 281701 29835
rect 281729 29807 281763 29835
rect 281791 29807 290577 29835
rect 290605 29807 290639 29835
rect 290667 29807 290701 29835
rect 290729 29807 290763 29835
rect 290791 29807 299256 29835
rect 299284 29807 299318 29835
rect 299346 29807 299380 29835
rect 299408 29807 299442 29835
rect 299470 29807 299998 29835
rect -6 29773 299998 29807
rect -6 29745 522 29773
rect 550 29745 584 29773
rect 612 29745 646 29773
rect 674 29745 708 29773
rect 736 29745 2577 29773
rect 2605 29745 2639 29773
rect 2667 29745 2701 29773
rect 2729 29745 2763 29773
rect 2791 29745 11577 29773
rect 11605 29745 11639 29773
rect 11667 29745 11701 29773
rect 11729 29745 11763 29773
rect 11791 29745 17259 29773
rect 17287 29745 17321 29773
rect 17349 29745 20577 29773
rect 20605 29745 20639 29773
rect 20667 29745 20701 29773
rect 20729 29745 20763 29773
rect 20791 29745 29577 29773
rect 29605 29745 29639 29773
rect 29667 29745 29701 29773
rect 29729 29745 29763 29773
rect 29791 29745 32619 29773
rect 32647 29745 32681 29773
rect 32709 29745 47979 29773
rect 48007 29745 48041 29773
rect 48069 29745 63339 29773
rect 63367 29745 63401 29773
rect 63429 29745 78699 29773
rect 78727 29745 78761 29773
rect 78789 29745 94059 29773
rect 94087 29745 94121 29773
rect 94149 29745 109419 29773
rect 109447 29745 109481 29773
rect 109509 29745 124779 29773
rect 124807 29745 124841 29773
rect 124869 29745 140139 29773
rect 140167 29745 140201 29773
rect 140229 29745 155499 29773
rect 155527 29745 155561 29773
rect 155589 29745 170859 29773
rect 170887 29745 170921 29773
rect 170949 29745 186219 29773
rect 186247 29745 186281 29773
rect 186309 29745 201579 29773
rect 201607 29745 201641 29773
rect 201669 29745 216939 29773
rect 216967 29745 217001 29773
rect 217029 29745 232299 29773
rect 232327 29745 232361 29773
rect 232389 29745 247659 29773
rect 247687 29745 247721 29773
rect 247749 29745 254577 29773
rect 254605 29745 254639 29773
rect 254667 29745 254701 29773
rect 254729 29745 254763 29773
rect 254791 29745 263577 29773
rect 263605 29745 263639 29773
rect 263667 29745 263701 29773
rect 263729 29745 263763 29773
rect 263791 29745 272577 29773
rect 272605 29745 272639 29773
rect 272667 29745 272701 29773
rect 272729 29745 272763 29773
rect 272791 29745 281577 29773
rect 281605 29745 281639 29773
rect 281667 29745 281701 29773
rect 281729 29745 281763 29773
rect 281791 29745 290577 29773
rect 290605 29745 290639 29773
rect 290667 29745 290701 29773
rect 290729 29745 290763 29773
rect 290791 29745 299256 29773
rect 299284 29745 299318 29773
rect 299346 29745 299380 29773
rect 299408 29745 299442 29773
rect 299470 29745 299998 29773
rect -6 29697 299998 29745
rect -6 23959 299998 24007
rect -6 23931 42 23959
rect 70 23931 104 23959
rect 132 23931 166 23959
rect 194 23931 228 23959
rect 256 23931 4437 23959
rect 4465 23931 4499 23959
rect 4527 23931 4561 23959
rect 4589 23931 4623 23959
rect 4651 23931 13437 23959
rect 13465 23931 13499 23959
rect 13527 23931 13561 23959
rect 13589 23931 13623 23959
rect 13651 23931 22437 23959
rect 22465 23931 22499 23959
rect 22527 23931 22561 23959
rect 22589 23931 22623 23959
rect 22651 23931 24939 23959
rect 24967 23931 25001 23959
rect 25029 23931 31437 23959
rect 31465 23931 31499 23959
rect 31527 23931 31561 23959
rect 31589 23931 31623 23959
rect 31651 23931 40299 23959
rect 40327 23931 40361 23959
rect 40389 23931 55659 23959
rect 55687 23931 55721 23959
rect 55749 23931 71019 23959
rect 71047 23931 71081 23959
rect 71109 23931 86379 23959
rect 86407 23931 86441 23959
rect 86469 23931 101739 23959
rect 101767 23931 101801 23959
rect 101829 23931 117099 23959
rect 117127 23931 117161 23959
rect 117189 23931 132459 23959
rect 132487 23931 132521 23959
rect 132549 23931 147819 23959
rect 147847 23931 147881 23959
rect 147909 23931 163179 23959
rect 163207 23931 163241 23959
rect 163269 23931 178539 23959
rect 178567 23931 178601 23959
rect 178629 23931 193899 23959
rect 193927 23931 193961 23959
rect 193989 23931 209259 23959
rect 209287 23931 209321 23959
rect 209349 23931 224619 23959
rect 224647 23931 224681 23959
rect 224709 23931 239979 23959
rect 240007 23931 240041 23959
rect 240069 23931 256437 23959
rect 256465 23931 256499 23959
rect 256527 23931 256561 23959
rect 256589 23931 256623 23959
rect 256651 23931 265437 23959
rect 265465 23931 265499 23959
rect 265527 23931 265561 23959
rect 265589 23931 265623 23959
rect 265651 23931 274437 23959
rect 274465 23931 274499 23959
rect 274527 23931 274561 23959
rect 274589 23931 274623 23959
rect 274651 23931 283437 23959
rect 283465 23931 283499 23959
rect 283527 23931 283561 23959
rect 283589 23931 283623 23959
rect 283651 23931 292437 23959
rect 292465 23931 292499 23959
rect 292527 23931 292561 23959
rect 292589 23931 292623 23959
rect 292651 23931 299736 23959
rect 299764 23931 299798 23959
rect 299826 23931 299860 23959
rect 299888 23931 299922 23959
rect 299950 23931 299998 23959
rect -6 23897 299998 23931
rect -6 23869 42 23897
rect 70 23869 104 23897
rect 132 23869 166 23897
rect 194 23869 228 23897
rect 256 23869 4437 23897
rect 4465 23869 4499 23897
rect 4527 23869 4561 23897
rect 4589 23869 4623 23897
rect 4651 23869 13437 23897
rect 13465 23869 13499 23897
rect 13527 23869 13561 23897
rect 13589 23869 13623 23897
rect 13651 23869 22437 23897
rect 22465 23869 22499 23897
rect 22527 23869 22561 23897
rect 22589 23869 22623 23897
rect 22651 23869 24939 23897
rect 24967 23869 25001 23897
rect 25029 23869 31437 23897
rect 31465 23869 31499 23897
rect 31527 23869 31561 23897
rect 31589 23869 31623 23897
rect 31651 23869 40299 23897
rect 40327 23869 40361 23897
rect 40389 23869 55659 23897
rect 55687 23869 55721 23897
rect 55749 23869 71019 23897
rect 71047 23869 71081 23897
rect 71109 23869 86379 23897
rect 86407 23869 86441 23897
rect 86469 23869 101739 23897
rect 101767 23869 101801 23897
rect 101829 23869 117099 23897
rect 117127 23869 117161 23897
rect 117189 23869 132459 23897
rect 132487 23869 132521 23897
rect 132549 23869 147819 23897
rect 147847 23869 147881 23897
rect 147909 23869 163179 23897
rect 163207 23869 163241 23897
rect 163269 23869 178539 23897
rect 178567 23869 178601 23897
rect 178629 23869 193899 23897
rect 193927 23869 193961 23897
rect 193989 23869 209259 23897
rect 209287 23869 209321 23897
rect 209349 23869 224619 23897
rect 224647 23869 224681 23897
rect 224709 23869 239979 23897
rect 240007 23869 240041 23897
rect 240069 23869 256437 23897
rect 256465 23869 256499 23897
rect 256527 23869 256561 23897
rect 256589 23869 256623 23897
rect 256651 23869 265437 23897
rect 265465 23869 265499 23897
rect 265527 23869 265561 23897
rect 265589 23869 265623 23897
rect 265651 23869 274437 23897
rect 274465 23869 274499 23897
rect 274527 23869 274561 23897
rect 274589 23869 274623 23897
rect 274651 23869 283437 23897
rect 283465 23869 283499 23897
rect 283527 23869 283561 23897
rect 283589 23869 283623 23897
rect 283651 23869 292437 23897
rect 292465 23869 292499 23897
rect 292527 23869 292561 23897
rect 292589 23869 292623 23897
rect 292651 23869 299736 23897
rect 299764 23869 299798 23897
rect 299826 23869 299860 23897
rect 299888 23869 299922 23897
rect 299950 23869 299998 23897
rect -6 23835 299998 23869
rect -6 23807 42 23835
rect 70 23807 104 23835
rect 132 23807 166 23835
rect 194 23807 228 23835
rect 256 23807 4437 23835
rect 4465 23807 4499 23835
rect 4527 23807 4561 23835
rect 4589 23807 4623 23835
rect 4651 23807 13437 23835
rect 13465 23807 13499 23835
rect 13527 23807 13561 23835
rect 13589 23807 13623 23835
rect 13651 23807 22437 23835
rect 22465 23807 22499 23835
rect 22527 23807 22561 23835
rect 22589 23807 22623 23835
rect 22651 23807 24939 23835
rect 24967 23807 25001 23835
rect 25029 23807 31437 23835
rect 31465 23807 31499 23835
rect 31527 23807 31561 23835
rect 31589 23807 31623 23835
rect 31651 23807 40299 23835
rect 40327 23807 40361 23835
rect 40389 23807 55659 23835
rect 55687 23807 55721 23835
rect 55749 23807 71019 23835
rect 71047 23807 71081 23835
rect 71109 23807 86379 23835
rect 86407 23807 86441 23835
rect 86469 23807 101739 23835
rect 101767 23807 101801 23835
rect 101829 23807 117099 23835
rect 117127 23807 117161 23835
rect 117189 23807 132459 23835
rect 132487 23807 132521 23835
rect 132549 23807 147819 23835
rect 147847 23807 147881 23835
rect 147909 23807 163179 23835
rect 163207 23807 163241 23835
rect 163269 23807 178539 23835
rect 178567 23807 178601 23835
rect 178629 23807 193899 23835
rect 193927 23807 193961 23835
rect 193989 23807 209259 23835
rect 209287 23807 209321 23835
rect 209349 23807 224619 23835
rect 224647 23807 224681 23835
rect 224709 23807 239979 23835
rect 240007 23807 240041 23835
rect 240069 23807 256437 23835
rect 256465 23807 256499 23835
rect 256527 23807 256561 23835
rect 256589 23807 256623 23835
rect 256651 23807 265437 23835
rect 265465 23807 265499 23835
rect 265527 23807 265561 23835
rect 265589 23807 265623 23835
rect 265651 23807 274437 23835
rect 274465 23807 274499 23835
rect 274527 23807 274561 23835
rect 274589 23807 274623 23835
rect 274651 23807 283437 23835
rect 283465 23807 283499 23835
rect 283527 23807 283561 23835
rect 283589 23807 283623 23835
rect 283651 23807 292437 23835
rect 292465 23807 292499 23835
rect 292527 23807 292561 23835
rect 292589 23807 292623 23835
rect 292651 23807 299736 23835
rect 299764 23807 299798 23835
rect 299826 23807 299860 23835
rect 299888 23807 299922 23835
rect 299950 23807 299998 23835
rect -6 23773 299998 23807
rect -6 23745 42 23773
rect 70 23745 104 23773
rect 132 23745 166 23773
rect 194 23745 228 23773
rect 256 23745 4437 23773
rect 4465 23745 4499 23773
rect 4527 23745 4561 23773
rect 4589 23745 4623 23773
rect 4651 23745 13437 23773
rect 13465 23745 13499 23773
rect 13527 23745 13561 23773
rect 13589 23745 13623 23773
rect 13651 23745 22437 23773
rect 22465 23745 22499 23773
rect 22527 23745 22561 23773
rect 22589 23745 22623 23773
rect 22651 23745 24939 23773
rect 24967 23745 25001 23773
rect 25029 23745 31437 23773
rect 31465 23745 31499 23773
rect 31527 23745 31561 23773
rect 31589 23745 31623 23773
rect 31651 23745 40299 23773
rect 40327 23745 40361 23773
rect 40389 23745 55659 23773
rect 55687 23745 55721 23773
rect 55749 23745 71019 23773
rect 71047 23745 71081 23773
rect 71109 23745 86379 23773
rect 86407 23745 86441 23773
rect 86469 23745 101739 23773
rect 101767 23745 101801 23773
rect 101829 23745 117099 23773
rect 117127 23745 117161 23773
rect 117189 23745 132459 23773
rect 132487 23745 132521 23773
rect 132549 23745 147819 23773
rect 147847 23745 147881 23773
rect 147909 23745 163179 23773
rect 163207 23745 163241 23773
rect 163269 23745 178539 23773
rect 178567 23745 178601 23773
rect 178629 23745 193899 23773
rect 193927 23745 193961 23773
rect 193989 23745 209259 23773
rect 209287 23745 209321 23773
rect 209349 23745 224619 23773
rect 224647 23745 224681 23773
rect 224709 23745 239979 23773
rect 240007 23745 240041 23773
rect 240069 23745 256437 23773
rect 256465 23745 256499 23773
rect 256527 23745 256561 23773
rect 256589 23745 256623 23773
rect 256651 23745 265437 23773
rect 265465 23745 265499 23773
rect 265527 23745 265561 23773
rect 265589 23745 265623 23773
rect 265651 23745 274437 23773
rect 274465 23745 274499 23773
rect 274527 23745 274561 23773
rect 274589 23745 274623 23773
rect 274651 23745 283437 23773
rect 283465 23745 283499 23773
rect 283527 23745 283561 23773
rect 283589 23745 283623 23773
rect 283651 23745 292437 23773
rect 292465 23745 292499 23773
rect 292527 23745 292561 23773
rect 292589 23745 292623 23773
rect 292651 23745 299736 23773
rect 299764 23745 299798 23773
rect 299826 23745 299860 23773
rect 299888 23745 299922 23773
rect 299950 23745 299998 23773
rect -6 23697 299998 23745
rect -6 20959 299998 21007
rect -6 20931 522 20959
rect 550 20931 584 20959
rect 612 20931 646 20959
rect 674 20931 708 20959
rect 736 20931 2577 20959
rect 2605 20931 2639 20959
rect 2667 20931 2701 20959
rect 2729 20931 2763 20959
rect 2791 20931 11577 20959
rect 11605 20931 11639 20959
rect 11667 20931 11701 20959
rect 11729 20931 11763 20959
rect 11791 20931 17259 20959
rect 17287 20931 17321 20959
rect 17349 20931 20577 20959
rect 20605 20931 20639 20959
rect 20667 20931 20701 20959
rect 20729 20931 20763 20959
rect 20791 20931 29577 20959
rect 29605 20931 29639 20959
rect 29667 20931 29701 20959
rect 29729 20931 29763 20959
rect 29791 20931 32619 20959
rect 32647 20931 32681 20959
rect 32709 20931 47979 20959
rect 48007 20931 48041 20959
rect 48069 20931 63339 20959
rect 63367 20931 63401 20959
rect 63429 20931 78699 20959
rect 78727 20931 78761 20959
rect 78789 20931 94059 20959
rect 94087 20931 94121 20959
rect 94149 20931 109419 20959
rect 109447 20931 109481 20959
rect 109509 20931 124779 20959
rect 124807 20931 124841 20959
rect 124869 20931 140139 20959
rect 140167 20931 140201 20959
rect 140229 20931 155499 20959
rect 155527 20931 155561 20959
rect 155589 20931 170859 20959
rect 170887 20931 170921 20959
rect 170949 20931 186219 20959
rect 186247 20931 186281 20959
rect 186309 20931 201579 20959
rect 201607 20931 201641 20959
rect 201669 20931 216939 20959
rect 216967 20931 217001 20959
rect 217029 20931 232299 20959
rect 232327 20931 232361 20959
rect 232389 20931 247659 20959
rect 247687 20931 247721 20959
rect 247749 20931 254577 20959
rect 254605 20931 254639 20959
rect 254667 20931 254701 20959
rect 254729 20931 254763 20959
rect 254791 20931 263577 20959
rect 263605 20931 263639 20959
rect 263667 20931 263701 20959
rect 263729 20931 263763 20959
rect 263791 20931 272577 20959
rect 272605 20931 272639 20959
rect 272667 20931 272701 20959
rect 272729 20931 272763 20959
rect 272791 20931 281577 20959
rect 281605 20931 281639 20959
rect 281667 20931 281701 20959
rect 281729 20931 281763 20959
rect 281791 20931 290577 20959
rect 290605 20931 290639 20959
rect 290667 20931 290701 20959
rect 290729 20931 290763 20959
rect 290791 20931 299256 20959
rect 299284 20931 299318 20959
rect 299346 20931 299380 20959
rect 299408 20931 299442 20959
rect 299470 20931 299998 20959
rect -6 20897 299998 20931
rect -6 20869 522 20897
rect 550 20869 584 20897
rect 612 20869 646 20897
rect 674 20869 708 20897
rect 736 20869 2577 20897
rect 2605 20869 2639 20897
rect 2667 20869 2701 20897
rect 2729 20869 2763 20897
rect 2791 20869 11577 20897
rect 11605 20869 11639 20897
rect 11667 20869 11701 20897
rect 11729 20869 11763 20897
rect 11791 20869 17259 20897
rect 17287 20869 17321 20897
rect 17349 20869 20577 20897
rect 20605 20869 20639 20897
rect 20667 20869 20701 20897
rect 20729 20869 20763 20897
rect 20791 20869 29577 20897
rect 29605 20869 29639 20897
rect 29667 20869 29701 20897
rect 29729 20869 29763 20897
rect 29791 20869 32619 20897
rect 32647 20869 32681 20897
rect 32709 20869 47979 20897
rect 48007 20869 48041 20897
rect 48069 20869 63339 20897
rect 63367 20869 63401 20897
rect 63429 20869 78699 20897
rect 78727 20869 78761 20897
rect 78789 20869 94059 20897
rect 94087 20869 94121 20897
rect 94149 20869 109419 20897
rect 109447 20869 109481 20897
rect 109509 20869 124779 20897
rect 124807 20869 124841 20897
rect 124869 20869 140139 20897
rect 140167 20869 140201 20897
rect 140229 20869 155499 20897
rect 155527 20869 155561 20897
rect 155589 20869 170859 20897
rect 170887 20869 170921 20897
rect 170949 20869 186219 20897
rect 186247 20869 186281 20897
rect 186309 20869 201579 20897
rect 201607 20869 201641 20897
rect 201669 20869 216939 20897
rect 216967 20869 217001 20897
rect 217029 20869 232299 20897
rect 232327 20869 232361 20897
rect 232389 20869 247659 20897
rect 247687 20869 247721 20897
rect 247749 20869 254577 20897
rect 254605 20869 254639 20897
rect 254667 20869 254701 20897
rect 254729 20869 254763 20897
rect 254791 20869 263577 20897
rect 263605 20869 263639 20897
rect 263667 20869 263701 20897
rect 263729 20869 263763 20897
rect 263791 20869 272577 20897
rect 272605 20869 272639 20897
rect 272667 20869 272701 20897
rect 272729 20869 272763 20897
rect 272791 20869 281577 20897
rect 281605 20869 281639 20897
rect 281667 20869 281701 20897
rect 281729 20869 281763 20897
rect 281791 20869 290577 20897
rect 290605 20869 290639 20897
rect 290667 20869 290701 20897
rect 290729 20869 290763 20897
rect 290791 20869 299256 20897
rect 299284 20869 299318 20897
rect 299346 20869 299380 20897
rect 299408 20869 299442 20897
rect 299470 20869 299998 20897
rect -6 20835 299998 20869
rect -6 20807 522 20835
rect 550 20807 584 20835
rect 612 20807 646 20835
rect 674 20807 708 20835
rect 736 20807 2577 20835
rect 2605 20807 2639 20835
rect 2667 20807 2701 20835
rect 2729 20807 2763 20835
rect 2791 20807 11577 20835
rect 11605 20807 11639 20835
rect 11667 20807 11701 20835
rect 11729 20807 11763 20835
rect 11791 20807 17259 20835
rect 17287 20807 17321 20835
rect 17349 20807 20577 20835
rect 20605 20807 20639 20835
rect 20667 20807 20701 20835
rect 20729 20807 20763 20835
rect 20791 20807 29577 20835
rect 29605 20807 29639 20835
rect 29667 20807 29701 20835
rect 29729 20807 29763 20835
rect 29791 20807 32619 20835
rect 32647 20807 32681 20835
rect 32709 20807 47979 20835
rect 48007 20807 48041 20835
rect 48069 20807 63339 20835
rect 63367 20807 63401 20835
rect 63429 20807 78699 20835
rect 78727 20807 78761 20835
rect 78789 20807 94059 20835
rect 94087 20807 94121 20835
rect 94149 20807 109419 20835
rect 109447 20807 109481 20835
rect 109509 20807 124779 20835
rect 124807 20807 124841 20835
rect 124869 20807 140139 20835
rect 140167 20807 140201 20835
rect 140229 20807 155499 20835
rect 155527 20807 155561 20835
rect 155589 20807 170859 20835
rect 170887 20807 170921 20835
rect 170949 20807 186219 20835
rect 186247 20807 186281 20835
rect 186309 20807 201579 20835
rect 201607 20807 201641 20835
rect 201669 20807 216939 20835
rect 216967 20807 217001 20835
rect 217029 20807 232299 20835
rect 232327 20807 232361 20835
rect 232389 20807 247659 20835
rect 247687 20807 247721 20835
rect 247749 20807 254577 20835
rect 254605 20807 254639 20835
rect 254667 20807 254701 20835
rect 254729 20807 254763 20835
rect 254791 20807 263577 20835
rect 263605 20807 263639 20835
rect 263667 20807 263701 20835
rect 263729 20807 263763 20835
rect 263791 20807 272577 20835
rect 272605 20807 272639 20835
rect 272667 20807 272701 20835
rect 272729 20807 272763 20835
rect 272791 20807 281577 20835
rect 281605 20807 281639 20835
rect 281667 20807 281701 20835
rect 281729 20807 281763 20835
rect 281791 20807 290577 20835
rect 290605 20807 290639 20835
rect 290667 20807 290701 20835
rect 290729 20807 290763 20835
rect 290791 20807 299256 20835
rect 299284 20807 299318 20835
rect 299346 20807 299380 20835
rect 299408 20807 299442 20835
rect 299470 20807 299998 20835
rect -6 20773 299998 20807
rect -6 20745 522 20773
rect 550 20745 584 20773
rect 612 20745 646 20773
rect 674 20745 708 20773
rect 736 20745 2577 20773
rect 2605 20745 2639 20773
rect 2667 20745 2701 20773
rect 2729 20745 2763 20773
rect 2791 20745 11577 20773
rect 11605 20745 11639 20773
rect 11667 20745 11701 20773
rect 11729 20745 11763 20773
rect 11791 20745 17259 20773
rect 17287 20745 17321 20773
rect 17349 20745 20577 20773
rect 20605 20745 20639 20773
rect 20667 20745 20701 20773
rect 20729 20745 20763 20773
rect 20791 20745 29577 20773
rect 29605 20745 29639 20773
rect 29667 20745 29701 20773
rect 29729 20745 29763 20773
rect 29791 20745 32619 20773
rect 32647 20745 32681 20773
rect 32709 20745 47979 20773
rect 48007 20745 48041 20773
rect 48069 20745 63339 20773
rect 63367 20745 63401 20773
rect 63429 20745 78699 20773
rect 78727 20745 78761 20773
rect 78789 20745 94059 20773
rect 94087 20745 94121 20773
rect 94149 20745 109419 20773
rect 109447 20745 109481 20773
rect 109509 20745 124779 20773
rect 124807 20745 124841 20773
rect 124869 20745 140139 20773
rect 140167 20745 140201 20773
rect 140229 20745 155499 20773
rect 155527 20745 155561 20773
rect 155589 20745 170859 20773
rect 170887 20745 170921 20773
rect 170949 20745 186219 20773
rect 186247 20745 186281 20773
rect 186309 20745 201579 20773
rect 201607 20745 201641 20773
rect 201669 20745 216939 20773
rect 216967 20745 217001 20773
rect 217029 20745 232299 20773
rect 232327 20745 232361 20773
rect 232389 20745 247659 20773
rect 247687 20745 247721 20773
rect 247749 20745 254577 20773
rect 254605 20745 254639 20773
rect 254667 20745 254701 20773
rect 254729 20745 254763 20773
rect 254791 20745 263577 20773
rect 263605 20745 263639 20773
rect 263667 20745 263701 20773
rect 263729 20745 263763 20773
rect 263791 20745 272577 20773
rect 272605 20745 272639 20773
rect 272667 20745 272701 20773
rect 272729 20745 272763 20773
rect 272791 20745 281577 20773
rect 281605 20745 281639 20773
rect 281667 20745 281701 20773
rect 281729 20745 281763 20773
rect 281791 20745 290577 20773
rect 290605 20745 290639 20773
rect 290667 20745 290701 20773
rect 290729 20745 290763 20773
rect 290791 20745 299256 20773
rect 299284 20745 299318 20773
rect 299346 20745 299380 20773
rect 299408 20745 299442 20773
rect 299470 20745 299998 20773
rect -6 20697 299998 20745
rect -6 14959 299998 15007
rect -6 14931 42 14959
rect 70 14931 104 14959
rect 132 14931 166 14959
rect 194 14931 228 14959
rect 256 14931 4437 14959
rect 4465 14931 4499 14959
rect 4527 14931 4561 14959
rect 4589 14931 4623 14959
rect 4651 14931 13437 14959
rect 13465 14931 13499 14959
rect 13527 14931 13561 14959
rect 13589 14931 13623 14959
rect 13651 14931 22437 14959
rect 22465 14931 22499 14959
rect 22527 14931 22561 14959
rect 22589 14931 22623 14959
rect 22651 14931 31437 14959
rect 31465 14931 31499 14959
rect 31527 14931 31561 14959
rect 31589 14931 31623 14959
rect 31651 14931 247437 14959
rect 247465 14931 247499 14959
rect 247527 14931 247561 14959
rect 247589 14931 247623 14959
rect 247651 14931 256437 14959
rect 256465 14931 256499 14959
rect 256527 14931 256561 14959
rect 256589 14931 256623 14959
rect 256651 14931 265437 14959
rect 265465 14931 265499 14959
rect 265527 14931 265561 14959
rect 265589 14931 265623 14959
rect 265651 14931 274437 14959
rect 274465 14931 274499 14959
rect 274527 14931 274561 14959
rect 274589 14931 274623 14959
rect 274651 14931 283437 14959
rect 283465 14931 283499 14959
rect 283527 14931 283561 14959
rect 283589 14931 283623 14959
rect 283651 14931 292437 14959
rect 292465 14931 292499 14959
rect 292527 14931 292561 14959
rect 292589 14931 292623 14959
rect 292651 14931 299736 14959
rect 299764 14931 299798 14959
rect 299826 14931 299860 14959
rect 299888 14931 299922 14959
rect 299950 14931 299998 14959
rect -6 14897 299998 14931
rect -6 14869 42 14897
rect 70 14869 104 14897
rect 132 14869 166 14897
rect 194 14869 228 14897
rect 256 14869 4437 14897
rect 4465 14869 4499 14897
rect 4527 14869 4561 14897
rect 4589 14869 4623 14897
rect 4651 14869 13437 14897
rect 13465 14869 13499 14897
rect 13527 14869 13561 14897
rect 13589 14869 13623 14897
rect 13651 14869 22437 14897
rect 22465 14869 22499 14897
rect 22527 14869 22561 14897
rect 22589 14869 22623 14897
rect 22651 14869 31437 14897
rect 31465 14869 31499 14897
rect 31527 14869 31561 14897
rect 31589 14869 31623 14897
rect 31651 14869 247437 14897
rect 247465 14869 247499 14897
rect 247527 14869 247561 14897
rect 247589 14869 247623 14897
rect 247651 14869 256437 14897
rect 256465 14869 256499 14897
rect 256527 14869 256561 14897
rect 256589 14869 256623 14897
rect 256651 14869 265437 14897
rect 265465 14869 265499 14897
rect 265527 14869 265561 14897
rect 265589 14869 265623 14897
rect 265651 14869 274437 14897
rect 274465 14869 274499 14897
rect 274527 14869 274561 14897
rect 274589 14869 274623 14897
rect 274651 14869 283437 14897
rect 283465 14869 283499 14897
rect 283527 14869 283561 14897
rect 283589 14869 283623 14897
rect 283651 14869 292437 14897
rect 292465 14869 292499 14897
rect 292527 14869 292561 14897
rect 292589 14869 292623 14897
rect 292651 14869 299736 14897
rect 299764 14869 299798 14897
rect 299826 14869 299860 14897
rect 299888 14869 299922 14897
rect 299950 14869 299998 14897
rect -6 14835 299998 14869
rect -6 14807 42 14835
rect 70 14807 104 14835
rect 132 14807 166 14835
rect 194 14807 228 14835
rect 256 14807 4437 14835
rect 4465 14807 4499 14835
rect 4527 14807 4561 14835
rect 4589 14807 4623 14835
rect 4651 14807 13437 14835
rect 13465 14807 13499 14835
rect 13527 14807 13561 14835
rect 13589 14807 13623 14835
rect 13651 14807 22437 14835
rect 22465 14807 22499 14835
rect 22527 14807 22561 14835
rect 22589 14807 22623 14835
rect 22651 14807 31437 14835
rect 31465 14807 31499 14835
rect 31527 14807 31561 14835
rect 31589 14807 31623 14835
rect 31651 14807 247437 14835
rect 247465 14807 247499 14835
rect 247527 14807 247561 14835
rect 247589 14807 247623 14835
rect 247651 14807 256437 14835
rect 256465 14807 256499 14835
rect 256527 14807 256561 14835
rect 256589 14807 256623 14835
rect 256651 14807 265437 14835
rect 265465 14807 265499 14835
rect 265527 14807 265561 14835
rect 265589 14807 265623 14835
rect 265651 14807 274437 14835
rect 274465 14807 274499 14835
rect 274527 14807 274561 14835
rect 274589 14807 274623 14835
rect 274651 14807 283437 14835
rect 283465 14807 283499 14835
rect 283527 14807 283561 14835
rect 283589 14807 283623 14835
rect 283651 14807 292437 14835
rect 292465 14807 292499 14835
rect 292527 14807 292561 14835
rect 292589 14807 292623 14835
rect 292651 14807 299736 14835
rect 299764 14807 299798 14835
rect 299826 14807 299860 14835
rect 299888 14807 299922 14835
rect 299950 14807 299998 14835
rect -6 14773 299998 14807
rect -6 14745 42 14773
rect 70 14745 104 14773
rect 132 14745 166 14773
rect 194 14745 228 14773
rect 256 14745 4437 14773
rect 4465 14745 4499 14773
rect 4527 14745 4561 14773
rect 4589 14745 4623 14773
rect 4651 14745 13437 14773
rect 13465 14745 13499 14773
rect 13527 14745 13561 14773
rect 13589 14745 13623 14773
rect 13651 14745 22437 14773
rect 22465 14745 22499 14773
rect 22527 14745 22561 14773
rect 22589 14745 22623 14773
rect 22651 14745 31437 14773
rect 31465 14745 31499 14773
rect 31527 14745 31561 14773
rect 31589 14745 31623 14773
rect 31651 14745 247437 14773
rect 247465 14745 247499 14773
rect 247527 14745 247561 14773
rect 247589 14745 247623 14773
rect 247651 14745 256437 14773
rect 256465 14745 256499 14773
rect 256527 14745 256561 14773
rect 256589 14745 256623 14773
rect 256651 14745 265437 14773
rect 265465 14745 265499 14773
rect 265527 14745 265561 14773
rect 265589 14745 265623 14773
rect 265651 14745 274437 14773
rect 274465 14745 274499 14773
rect 274527 14745 274561 14773
rect 274589 14745 274623 14773
rect 274651 14745 283437 14773
rect 283465 14745 283499 14773
rect 283527 14745 283561 14773
rect 283589 14745 283623 14773
rect 283651 14745 292437 14773
rect 292465 14745 292499 14773
rect 292527 14745 292561 14773
rect 292589 14745 292623 14773
rect 292651 14745 299736 14773
rect 299764 14745 299798 14773
rect 299826 14745 299860 14773
rect 299888 14745 299922 14773
rect 299950 14745 299998 14773
rect -6 14697 299998 14745
rect -6 11959 299998 12007
rect -6 11931 522 11959
rect 550 11931 584 11959
rect 612 11931 646 11959
rect 674 11931 708 11959
rect 736 11931 2577 11959
rect 2605 11931 2639 11959
rect 2667 11931 2701 11959
rect 2729 11931 2763 11959
rect 2791 11931 11577 11959
rect 11605 11931 11639 11959
rect 11667 11931 11701 11959
rect 11729 11931 11763 11959
rect 11791 11931 20577 11959
rect 20605 11931 20639 11959
rect 20667 11931 20701 11959
rect 20729 11931 20763 11959
rect 20791 11931 29577 11959
rect 29605 11931 29639 11959
rect 29667 11931 29701 11959
rect 29729 11931 29763 11959
rect 29791 11931 38577 11959
rect 38605 11931 38639 11959
rect 38667 11931 38701 11959
rect 38729 11931 38763 11959
rect 38791 11931 47577 11959
rect 47605 11931 47639 11959
rect 47667 11931 47701 11959
rect 47729 11931 47763 11959
rect 47791 11931 56577 11959
rect 56605 11931 56639 11959
rect 56667 11931 56701 11959
rect 56729 11931 56763 11959
rect 56791 11931 65577 11959
rect 65605 11931 65639 11959
rect 65667 11931 65701 11959
rect 65729 11931 65763 11959
rect 65791 11931 74577 11959
rect 74605 11931 74639 11959
rect 74667 11931 74701 11959
rect 74729 11931 74763 11959
rect 74791 11931 83577 11959
rect 83605 11931 83639 11959
rect 83667 11931 83701 11959
rect 83729 11931 83763 11959
rect 83791 11931 92577 11959
rect 92605 11931 92639 11959
rect 92667 11931 92701 11959
rect 92729 11931 92763 11959
rect 92791 11931 101577 11959
rect 101605 11931 101639 11959
rect 101667 11931 101701 11959
rect 101729 11931 101763 11959
rect 101791 11931 110577 11959
rect 110605 11931 110639 11959
rect 110667 11931 110701 11959
rect 110729 11931 110763 11959
rect 110791 11931 119577 11959
rect 119605 11931 119639 11959
rect 119667 11931 119701 11959
rect 119729 11931 119763 11959
rect 119791 11931 128577 11959
rect 128605 11931 128639 11959
rect 128667 11931 128701 11959
rect 128729 11931 128763 11959
rect 128791 11931 137577 11959
rect 137605 11931 137639 11959
rect 137667 11931 137701 11959
rect 137729 11931 137763 11959
rect 137791 11931 146577 11959
rect 146605 11931 146639 11959
rect 146667 11931 146701 11959
rect 146729 11931 146763 11959
rect 146791 11931 155577 11959
rect 155605 11931 155639 11959
rect 155667 11931 155701 11959
rect 155729 11931 155763 11959
rect 155791 11931 164577 11959
rect 164605 11931 164639 11959
rect 164667 11931 164701 11959
rect 164729 11931 164763 11959
rect 164791 11931 173577 11959
rect 173605 11931 173639 11959
rect 173667 11931 173701 11959
rect 173729 11931 173763 11959
rect 173791 11931 182577 11959
rect 182605 11931 182639 11959
rect 182667 11931 182701 11959
rect 182729 11931 182763 11959
rect 182791 11931 191577 11959
rect 191605 11931 191639 11959
rect 191667 11931 191701 11959
rect 191729 11931 191763 11959
rect 191791 11931 200577 11959
rect 200605 11931 200639 11959
rect 200667 11931 200701 11959
rect 200729 11931 200763 11959
rect 200791 11931 209577 11959
rect 209605 11931 209639 11959
rect 209667 11931 209701 11959
rect 209729 11931 209763 11959
rect 209791 11931 218577 11959
rect 218605 11931 218639 11959
rect 218667 11931 218701 11959
rect 218729 11931 218763 11959
rect 218791 11931 227577 11959
rect 227605 11931 227639 11959
rect 227667 11931 227701 11959
rect 227729 11931 227763 11959
rect 227791 11931 236577 11959
rect 236605 11931 236639 11959
rect 236667 11931 236701 11959
rect 236729 11931 236763 11959
rect 236791 11931 245577 11959
rect 245605 11931 245639 11959
rect 245667 11931 245701 11959
rect 245729 11931 245763 11959
rect 245791 11931 254577 11959
rect 254605 11931 254639 11959
rect 254667 11931 254701 11959
rect 254729 11931 254763 11959
rect 254791 11931 263577 11959
rect 263605 11931 263639 11959
rect 263667 11931 263701 11959
rect 263729 11931 263763 11959
rect 263791 11931 272577 11959
rect 272605 11931 272639 11959
rect 272667 11931 272701 11959
rect 272729 11931 272763 11959
rect 272791 11931 281577 11959
rect 281605 11931 281639 11959
rect 281667 11931 281701 11959
rect 281729 11931 281763 11959
rect 281791 11931 290577 11959
rect 290605 11931 290639 11959
rect 290667 11931 290701 11959
rect 290729 11931 290763 11959
rect 290791 11931 299256 11959
rect 299284 11931 299318 11959
rect 299346 11931 299380 11959
rect 299408 11931 299442 11959
rect 299470 11931 299998 11959
rect -6 11897 299998 11931
rect -6 11869 522 11897
rect 550 11869 584 11897
rect 612 11869 646 11897
rect 674 11869 708 11897
rect 736 11869 2577 11897
rect 2605 11869 2639 11897
rect 2667 11869 2701 11897
rect 2729 11869 2763 11897
rect 2791 11869 11577 11897
rect 11605 11869 11639 11897
rect 11667 11869 11701 11897
rect 11729 11869 11763 11897
rect 11791 11869 20577 11897
rect 20605 11869 20639 11897
rect 20667 11869 20701 11897
rect 20729 11869 20763 11897
rect 20791 11869 29577 11897
rect 29605 11869 29639 11897
rect 29667 11869 29701 11897
rect 29729 11869 29763 11897
rect 29791 11869 38577 11897
rect 38605 11869 38639 11897
rect 38667 11869 38701 11897
rect 38729 11869 38763 11897
rect 38791 11869 47577 11897
rect 47605 11869 47639 11897
rect 47667 11869 47701 11897
rect 47729 11869 47763 11897
rect 47791 11869 56577 11897
rect 56605 11869 56639 11897
rect 56667 11869 56701 11897
rect 56729 11869 56763 11897
rect 56791 11869 65577 11897
rect 65605 11869 65639 11897
rect 65667 11869 65701 11897
rect 65729 11869 65763 11897
rect 65791 11869 74577 11897
rect 74605 11869 74639 11897
rect 74667 11869 74701 11897
rect 74729 11869 74763 11897
rect 74791 11869 83577 11897
rect 83605 11869 83639 11897
rect 83667 11869 83701 11897
rect 83729 11869 83763 11897
rect 83791 11869 92577 11897
rect 92605 11869 92639 11897
rect 92667 11869 92701 11897
rect 92729 11869 92763 11897
rect 92791 11869 101577 11897
rect 101605 11869 101639 11897
rect 101667 11869 101701 11897
rect 101729 11869 101763 11897
rect 101791 11869 110577 11897
rect 110605 11869 110639 11897
rect 110667 11869 110701 11897
rect 110729 11869 110763 11897
rect 110791 11869 119577 11897
rect 119605 11869 119639 11897
rect 119667 11869 119701 11897
rect 119729 11869 119763 11897
rect 119791 11869 128577 11897
rect 128605 11869 128639 11897
rect 128667 11869 128701 11897
rect 128729 11869 128763 11897
rect 128791 11869 137577 11897
rect 137605 11869 137639 11897
rect 137667 11869 137701 11897
rect 137729 11869 137763 11897
rect 137791 11869 146577 11897
rect 146605 11869 146639 11897
rect 146667 11869 146701 11897
rect 146729 11869 146763 11897
rect 146791 11869 155577 11897
rect 155605 11869 155639 11897
rect 155667 11869 155701 11897
rect 155729 11869 155763 11897
rect 155791 11869 164577 11897
rect 164605 11869 164639 11897
rect 164667 11869 164701 11897
rect 164729 11869 164763 11897
rect 164791 11869 173577 11897
rect 173605 11869 173639 11897
rect 173667 11869 173701 11897
rect 173729 11869 173763 11897
rect 173791 11869 182577 11897
rect 182605 11869 182639 11897
rect 182667 11869 182701 11897
rect 182729 11869 182763 11897
rect 182791 11869 191577 11897
rect 191605 11869 191639 11897
rect 191667 11869 191701 11897
rect 191729 11869 191763 11897
rect 191791 11869 200577 11897
rect 200605 11869 200639 11897
rect 200667 11869 200701 11897
rect 200729 11869 200763 11897
rect 200791 11869 209577 11897
rect 209605 11869 209639 11897
rect 209667 11869 209701 11897
rect 209729 11869 209763 11897
rect 209791 11869 218577 11897
rect 218605 11869 218639 11897
rect 218667 11869 218701 11897
rect 218729 11869 218763 11897
rect 218791 11869 227577 11897
rect 227605 11869 227639 11897
rect 227667 11869 227701 11897
rect 227729 11869 227763 11897
rect 227791 11869 236577 11897
rect 236605 11869 236639 11897
rect 236667 11869 236701 11897
rect 236729 11869 236763 11897
rect 236791 11869 245577 11897
rect 245605 11869 245639 11897
rect 245667 11869 245701 11897
rect 245729 11869 245763 11897
rect 245791 11869 254577 11897
rect 254605 11869 254639 11897
rect 254667 11869 254701 11897
rect 254729 11869 254763 11897
rect 254791 11869 263577 11897
rect 263605 11869 263639 11897
rect 263667 11869 263701 11897
rect 263729 11869 263763 11897
rect 263791 11869 272577 11897
rect 272605 11869 272639 11897
rect 272667 11869 272701 11897
rect 272729 11869 272763 11897
rect 272791 11869 281577 11897
rect 281605 11869 281639 11897
rect 281667 11869 281701 11897
rect 281729 11869 281763 11897
rect 281791 11869 290577 11897
rect 290605 11869 290639 11897
rect 290667 11869 290701 11897
rect 290729 11869 290763 11897
rect 290791 11869 299256 11897
rect 299284 11869 299318 11897
rect 299346 11869 299380 11897
rect 299408 11869 299442 11897
rect 299470 11869 299998 11897
rect -6 11835 299998 11869
rect -6 11807 522 11835
rect 550 11807 584 11835
rect 612 11807 646 11835
rect 674 11807 708 11835
rect 736 11807 2577 11835
rect 2605 11807 2639 11835
rect 2667 11807 2701 11835
rect 2729 11807 2763 11835
rect 2791 11807 11577 11835
rect 11605 11807 11639 11835
rect 11667 11807 11701 11835
rect 11729 11807 11763 11835
rect 11791 11807 20577 11835
rect 20605 11807 20639 11835
rect 20667 11807 20701 11835
rect 20729 11807 20763 11835
rect 20791 11807 29577 11835
rect 29605 11807 29639 11835
rect 29667 11807 29701 11835
rect 29729 11807 29763 11835
rect 29791 11807 38577 11835
rect 38605 11807 38639 11835
rect 38667 11807 38701 11835
rect 38729 11807 38763 11835
rect 38791 11807 47577 11835
rect 47605 11807 47639 11835
rect 47667 11807 47701 11835
rect 47729 11807 47763 11835
rect 47791 11807 56577 11835
rect 56605 11807 56639 11835
rect 56667 11807 56701 11835
rect 56729 11807 56763 11835
rect 56791 11807 65577 11835
rect 65605 11807 65639 11835
rect 65667 11807 65701 11835
rect 65729 11807 65763 11835
rect 65791 11807 74577 11835
rect 74605 11807 74639 11835
rect 74667 11807 74701 11835
rect 74729 11807 74763 11835
rect 74791 11807 83577 11835
rect 83605 11807 83639 11835
rect 83667 11807 83701 11835
rect 83729 11807 83763 11835
rect 83791 11807 92577 11835
rect 92605 11807 92639 11835
rect 92667 11807 92701 11835
rect 92729 11807 92763 11835
rect 92791 11807 101577 11835
rect 101605 11807 101639 11835
rect 101667 11807 101701 11835
rect 101729 11807 101763 11835
rect 101791 11807 110577 11835
rect 110605 11807 110639 11835
rect 110667 11807 110701 11835
rect 110729 11807 110763 11835
rect 110791 11807 119577 11835
rect 119605 11807 119639 11835
rect 119667 11807 119701 11835
rect 119729 11807 119763 11835
rect 119791 11807 128577 11835
rect 128605 11807 128639 11835
rect 128667 11807 128701 11835
rect 128729 11807 128763 11835
rect 128791 11807 137577 11835
rect 137605 11807 137639 11835
rect 137667 11807 137701 11835
rect 137729 11807 137763 11835
rect 137791 11807 146577 11835
rect 146605 11807 146639 11835
rect 146667 11807 146701 11835
rect 146729 11807 146763 11835
rect 146791 11807 155577 11835
rect 155605 11807 155639 11835
rect 155667 11807 155701 11835
rect 155729 11807 155763 11835
rect 155791 11807 164577 11835
rect 164605 11807 164639 11835
rect 164667 11807 164701 11835
rect 164729 11807 164763 11835
rect 164791 11807 173577 11835
rect 173605 11807 173639 11835
rect 173667 11807 173701 11835
rect 173729 11807 173763 11835
rect 173791 11807 182577 11835
rect 182605 11807 182639 11835
rect 182667 11807 182701 11835
rect 182729 11807 182763 11835
rect 182791 11807 191577 11835
rect 191605 11807 191639 11835
rect 191667 11807 191701 11835
rect 191729 11807 191763 11835
rect 191791 11807 200577 11835
rect 200605 11807 200639 11835
rect 200667 11807 200701 11835
rect 200729 11807 200763 11835
rect 200791 11807 209577 11835
rect 209605 11807 209639 11835
rect 209667 11807 209701 11835
rect 209729 11807 209763 11835
rect 209791 11807 218577 11835
rect 218605 11807 218639 11835
rect 218667 11807 218701 11835
rect 218729 11807 218763 11835
rect 218791 11807 227577 11835
rect 227605 11807 227639 11835
rect 227667 11807 227701 11835
rect 227729 11807 227763 11835
rect 227791 11807 236577 11835
rect 236605 11807 236639 11835
rect 236667 11807 236701 11835
rect 236729 11807 236763 11835
rect 236791 11807 245577 11835
rect 245605 11807 245639 11835
rect 245667 11807 245701 11835
rect 245729 11807 245763 11835
rect 245791 11807 254577 11835
rect 254605 11807 254639 11835
rect 254667 11807 254701 11835
rect 254729 11807 254763 11835
rect 254791 11807 263577 11835
rect 263605 11807 263639 11835
rect 263667 11807 263701 11835
rect 263729 11807 263763 11835
rect 263791 11807 272577 11835
rect 272605 11807 272639 11835
rect 272667 11807 272701 11835
rect 272729 11807 272763 11835
rect 272791 11807 281577 11835
rect 281605 11807 281639 11835
rect 281667 11807 281701 11835
rect 281729 11807 281763 11835
rect 281791 11807 290577 11835
rect 290605 11807 290639 11835
rect 290667 11807 290701 11835
rect 290729 11807 290763 11835
rect 290791 11807 299256 11835
rect 299284 11807 299318 11835
rect 299346 11807 299380 11835
rect 299408 11807 299442 11835
rect 299470 11807 299998 11835
rect -6 11773 299998 11807
rect -6 11745 522 11773
rect 550 11745 584 11773
rect 612 11745 646 11773
rect 674 11745 708 11773
rect 736 11745 2577 11773
rect 2605 11745 2639 11773
rect 2667 11745 2701 11773
rect 2729 11745 2763 11773
rect 2791 11745 11577 11773
rect 11605 11745 11639 11773
rect 11667 11745 11701 11773
rect 11729 11745 11763 11773
rect 11791 11745 20577 11773
rect 20605 11745 20639 11773
rect 20667 11745 20701 11773
rect 20729 11745 20763 11773
rect 20791 11745 29577 11773
rect 29605 11745 29639 11773
rect 29667 11745 29701 11773
rect 29729 11745 29763 11773
rect 29791 11745 38577 11773
rect 38605 11745 38639 11773
rect 38667 11745 38701 11773
rect 38729 11745 38763 11773
rect 38791 11745 47577 11773
rect 47605 11745 47639 11773
rect 47667 11745 47701 11773
rect 47729 11745 47763 11773
rect 47791 11745 56577 11773
rect 56605 11745 56639 11773
rect 56667 11745 56701 11773
rect 56729 11745 56763 11773
rect 56791 11745 65577 11773
rect 65605 11745 65639 11773
rect 65667 11745 65701 11773
rect 65729 11745 65763 11773
rect 65791 11745 74577 11773
rect 74605 11745 74639 11773
rect 74667 11745 74701 11773
rect 74729 11745 74763 11773
rect 74791 11745 83577 11773
rect 83605 11745 83639 11773
rect 83667 11745 83701 11773
rect 83729 11745 83763 11773
rect 83791 11745 92577 11773
rect 92605 11745 92639 11773
rect 92667 11745 92701 11773
rect 92729 11745 92763 11773
rect 92791 11745 101577 11773
rect 101605 11745 101639 11773
rect 101667 11745 101701 11773
rect 101729 11745 101763 11773
rect 101791 11745 110577 11773
rect 110605 11745 110639 11773
rect 110667 11745 110701 11773
rect 110729 11745 110763 11773
rect 110791 11745 119577 11773
rect 119605 11745 119639 11773
rect 119667 11745 119701 11773
rect 119729 11745 119763 11773
rect 119791 11745 128577 11773
rect 128605 11745 128639 11773
rect 128667 11745 128701 11773
rect 128729 11745 128763 11773
rect 128791 11745 137577 11773
rect 137605 11745 137639 11773
rect 137667 11745 137701 11773
rect 137729 11745 137763 11773
rect 137791 11745 146577 11773
rect 146605 11745 146639 11773
rect 146667 11745 146701 11773
rect 146729 11745 146763 11773
rect 146791 11745 155577 11773
rect 155605 11745 155639 11773
rect 155667 11745 155701 11773
rect 155729 11745 155763 11773
rect 155791 11745 164577 11773
rect 164605 11745 164639 11773
rect 164667 11745 164701 11773
rect 164729 11745 164763 11773
rect 164791 11745 173577 11773
rect 173605 11745 173639 11773
rect 173667 11745 173701 11773
rect 173729 11745 173763 11773
rect 173791 11745 182577 11773
rect 182605 11745 182639 11773
rect 182667 11745 182701 11773
rect 182729 11745 182763 11773
rect 182791 11745 191577 11773
rect 191605 11745 191639 11773
rect 191667 11745 191701 11773
rect 191729 11745 191763 11773
rect 191791 11745 200577 11773
rect 200605 11745 200639 11773
rect 200667 11745 200701 11773
rect 200729 11745 200763 11773
rect 200791 11745 209577 11773
rect 209605 11745 209639 11773
rect 209667 11745 209701 11773
rect 209729 11745 209763 11773
rect 209791 11745 218577 11773
rect 218605 11745 218639 11773
rect 218667 11745 218701 11773
rect 218729 11745 218763 11773
rect 218791 11745 227577 11773
rect 227605 11745 227639 11773
rect 227667 11745 227701 11773
rect 227729 11745 227763 11773
rect 227791 11745 236577 11773
rect 236605 11745 236639 11773
rect 236667 11745 236701 11773
rect 236729 11745 236763 11773
rect 236791 11745 245577 11773
rect 245605 11745 245639 11773
rect 245667 11745 245701 11773
rect 245729 11745 245763 11773
rect 245791 11745 254577 11773
rect 254605 11745 254639 11773
rect 254667 11745 254701 11773
rect 254729 11745 254763 11773
rect 254791 11745 263577 11773
rect 263605 11745 263639 11773
rect 263667 11745 263701 11773
rect 263729 11745 263763 11773
rect 263791 11745 272577 11773
rect 272605 11745 272639 11773
rect 272667 11745 272701 11773
rect 272729 11745 272763 11773
rect 272791 11745 281577 11773
rect 281605 11745 281639 11773
rect 281667 11745 281701 11773
rect 281729 11745 281763 11773
rect 281791 11745 290577 11773
rect 290605 11745 290639 11773
rect 290667 11745 290701 11773
rect 290729 11745 290763 11773
rect 290791 11745 299256 11773
rect 299284 11745 299318 11773
rect 299346 11745 299380 11773
rect 299408 11745 299442 11773
rect 299470 11745 299998 11773
rect -6 11697 299998 11745
rect -6 5959 299998 6007
rect -6 5931 42 5959
rect 70 5931 104 5959
rect 132 5931 166 5959
rect 194 5931 228 5959
rect 256 5931 4437 5959
rect 4465 5931 4499 5959
rect 4527 5931 4561 5959
rect 4589 5931 4623 5959
rect 4651 5931 13437 5959
rect 13465 5931 13499 5959
rect 13527 5931 13561 5959
rect 13589 5931 13623 5959
rect 13651 5931 22437 5959
rect 22465 5931 22499 5959
rect 22527 5931 22561 5959
rect 22589 5931 22623 5959
rect 22651 5931 31437 5959
rect 31465 5931 31499 5959
rect 31527 5931 31561 5959
rect 31589 5931 31623 5959
rect 31651 5931 40437 5959
rect 40465 5931 40499 5959
rect 40527 5931 40561 5959
rect 40589 5931 40623 5959
rect 40651 5931 49437 5959
rect 49465 5931 49499 5959
rect 49527 5931 49561 5959
rect 49589 5931 49623 5959
rect 49651 5931 58437 5959
rect 58465 5931 58499 5959
rect 58527 5931 58561 5959
rect 58589 5931 58623 5959
rect 58651 5931 67437 5959
rect 67465 5931 67499 5959
rect 67527 5931 67561 5959
rect 67589 5931 67623 5959
rect 67651 5931 76437 5959
rect 76465 5931 76499 5959
rect 76527 5931 76561 5959
rect 76589 5931 76623 5959
rect 76651 5931 85437 5959
rect 85465 5931 85499 5959
rect 85527 5931 85561 5959
rect 85589 5931 85623 5959
rect 85651 5931 94437 5959
rect 94465 5931 94499 5959
rect 94527 5931 94561 5959
rect 94589 5931 94623 5959
rect 94651 5931 103437 5959
rect 103465 5931 103499 5959
rect 103527 5931 103561 5959
rect 103589 5931 103623 5959
rect 103651 5931 112437 5959
rect 112465 5931 112499 5959
rect 112527 5931 112561 5959
rect 112589 5931 112623 5959
rect 112651 5931 121437 5959
rect 121465 5931 121499 5959
rect 121527 5931 121561 5959
rect 121589 5931 121623 5959
rect 121651 5931 130437 5959
rect 130465 5931 130499 5959
rect 130527 5931 130561 5959
rect 130589 5931 130623 5959
rect 130651 5931 139437 5959
rect 139465 5931 139499 5959
rect 139527 5931 139561 5959
rect 139589 5931 139623 5959
rect 139651 5931 148437 5959
rect 148465 5931 148499 5959
rect 148527 5931 148561 5959
rect 148589 5931 148623 5959
rect 148651 5931 157437 5959
rect 157465 5931 157499 5959
rect 157527 5931 157561 5959
rect 157589 5931 157623 5959
rect 157651 5931 166437 5959
rect 166465 5931 166499 5959
rect 166527 5931 166561 5959
rect 166589 5931 166623 5959
rect 166651 5931 175437 5959
rect 175465 5931 175499 5959
rect 175527 5931 175561 5959
rect 175589 5931 175623 5959
rect 175651 5931 184437 5959
rect 184465 5931 184499 5959
rect 184527 5931 184561 5959
rect 184589 5931 184623 5959
rect 184651 5931 193437 5959
rect 193465 5931 193499 5959
rect 193527 5931 193561 5959
rect 193589 5931 193623 5959
rect 193651 5931 202437 5959
rect 202465 5931 202499 5959
rect 202527 5931 202561 5959
rect 202589 5931 202623 5959
rect 202651 5931 211437 5959
rect 211465 5931 211499 5959
rect 211527 5931 211561 5959
rect 211589 5931 211623 5959
rect 211651 5931 220437 5959
rect 220465 5931 220499 5959
rect 220527 5931 220561 5959
rect 220589 5931 220623 5959
rect 220651 5931 229437 5959
rect 229465 5931 229499 5959
rect 229527 5931 229561 5959
rect 229589 5931 229623 5959
rect 229651 5931 238437 5959
rect 238465 5931 238499 5959
rect 238527 5931 238561 5959
rect 238589 5931 238623 5959
rect 238651 5931 247437 5959
rect 247465 5931 247499 5959
rect 247527 5931 247561 5959
rect 247589 5931 247623 5959
rect 247651 5931 256437 5959
rect 256465 5931 256499 5959
rect 256527 5931 256561 5959
rect 256589 5931 256623 5959
rect 256651 5931 265437 5959
rect 265465 5931 265499 5959
rect 265527 5931 265561 5959
rect 265589 5931 265623 5959
rect 265651 5931 274437 5959
rect 274465 5931 274499 5959
rect 274527 5931 274561 5959
rect 274589 5931 274623 5959
rect 274651 5931 283437 5959
rect 283465 5931 283499 5959
rect 283527 5931 283561 5959
rect 283589 5931 283623 5959
rect 283651 5931 292437 5959
rect 292465 5931 292499 5959
rect 292527 5931 292561 5959
rect 292589 5931 292623 5959
rect 292651 5931 299736 5959
rect 299764 5931 299798 5959
rect 299826 5931 299860 5959
rect 299888 5931 299922 5959
rect 299950 5931 299998 5959
rect -6 5897 299998 5931
rect -6 5869 42 5897
rect 70 5869 104 5897
rect 132 5869 166 5897
rect 194 5869 228 5897
rect 256 5869 4437 5897
rect 4465 5869 4499 5897
rect 4527 5869 4561 5897
rect 4589 5869 4623 5897
rect 4651 5869 13437 5897
rect 13465 5869 13499 5897
rect 13527 5869 13561 5897
rect 13589 5869 13623 5897
rect 13651 5869 22437 5897
rect 22465 5869 22499 5897
rect 22527 5869 22561 5897
rect 22589 5869 22623 5897
rect 22651 5869 31437 5897
rect 31465 5869 31499 5897
rect 31527 5869 31561 5897
rect 31589 5869 31623 5897
rect 31651 5869 40437 5897
rect 40465 5869 40499 5897
rect 40527 5869 40561 5897
rect 40589 5869 40623 5897
rect 40651 5869 49437 5897
rect 49465 5869 49499 5897
rect 49527 5869 49561 5897
rect 49589 5869 49623 5897
rect 49651 5869 58437 5897
rect 58465 5869 58499 5897
rect 58527 5869 58561 5897
rect 58589 5869 58623 5897
rect 58651 5869 67437 5897
rect 67465 5869 67499 5897
rect 67527 5869 67561 5897
rect 67589 5869 67623 5897
rect 67651 5869 76437 5897
rect 76465 5869 76499 5897
rect 76527 5869 76561 5897
rect 76589 5869 76623 5897
rect 76651 5869 85437 5897
rect 85465 5869 85499 5897
rect 85527 5869 85561 5897
rect 85589 5869 85623 5897
rect 85651 5869 94437 5897
rect 94465 5869 94499 5897
rect 94527 5869 94561 5897
rect 94589 5869 94623 5897
rect 94651 5869 103437 5897
rect 103465 5869 103499 5897
rect 103527 5869 103561 5897
rect 103589 5869 103623 5897
rect 103651 5869 112437 5897
rect 112465 5869 112499 5897
rect 112527 5869 112561 5897
rect 112589 5869 112623 5897
rect 112651 5869 121437 5897
rect 121465 5869 121499 5897
rect 121527 5869 121561 5897
rect 121589 5869 121623 5897
rect 121651 5869 130437 5897
rect 130465 5869 130499 5897
rect 130527 5869 130561 5897
rect 130589 5869 130623 5897
rect 130651 5869 139437 5897
rect 139465 5869 139499 5897
rect 139527 5869 139561 5897
rect 139589 5869 139623 5897
rect 139651 5869 148437 5897
rect 148465 5869 148499 5897
rect 148527 5869 148561 5897
rect 148589 5869 148623 5897
rect 148651 5869 157437 5897
rect 157465 5869 157499 5897
rect 157527 5869 157561 5897
rect 157589 5869 157623 5897
rect 157651 5869 166437 5897
rect 166465 5869 166499 5897
rect 166527 5869 166561 5897
rect 166589 5869 166623 5897
rect 166651 5869 175437 5897
rect 175465 5869 175499 5897
rect 175527 5869 175561 5897
rect 175589 5869 175623 5897
rect 175651 5869 184437 5897
rect 184465 5869 184499 5897
rect 184527 5869 184561 5897
rect 184589 5869 184623 5897
rect 184651 5869 193437 5897
rect 193465 5869 193499 5897
rect 193527 5869 193561 5897
rect 193589 5869 193623 5897
rect 193651 5869 202437 5897
rect 202465 5869 202499 5897
rect 202527 5869 202561 5897
rect 202589 5869 202623 5897
rect 202651 5869 211437 5897
rect 211465 5869 211499 5897
rect 211527 5869 211561 5897
rect 211589 5869 211623 5897
rect 211651 5869 220437 5897
rect 220465 5869 220499 5897
rect 220527 5869 220561 5897
rect 220589 5869 220623 5897
rect 220651 5869 229437 5897
rect 229465 5869 229499 5897
rect 229527 5869 229561 5897
rect 229589 5869 229623 5897
rect 229651 5869 238437 5897
rect 238465 5869 238499 5897
rect 238527 5869 238561 5897
rect 238589 5869 238623 5897
rect 238651 5869 247437 5897
rect 247465 5869 247499 5897
rect 247527 5869 247561 5897
rect 247589 5869 247623 5897
rect 247651 5869 256437 5897
rect 256465 5869 256499 5897
rect 256527 5869 256561 5897
rect 256589 5869 256623 5897
rect 256651 5869 265437 5897
rect 265465 5869 265499 5897
rect 265527 5869 265561 5897
rect 265589 5869 265623 5897
rect 265651 5869 274437 5897
rect 274465 5869 274499 5897
rect 274527 5869 274561 5897
rect 274589 5869 274623 5897
rect 274651 5869 283437 5897
rect 283465 5869 283499 5897
rect 283527 5869 283561 5897
rect 283589 5869 283623 5897
rect 283651 5869 292437 5897
rect 292465 5869 292499 5897
rect 292527 5869 292561 5897
rect 292589 5869 292623 5897
rect 292651 5869 299736 5897
rect 299764 5869 299798 5897
rect 299826 5869 299860 5897
rect 299888 5869 299922 5897
rect 299950 5869 299998 5897
rect -6 5835 299998 5869
rect -6 5807 42 5835
rect 70 5807 104 5835
rect 132 5807 166 5835
rect 194 5807 228 5835
rect 256 5807 4437 5835
rect 4465 5807 4499 5835
rect 4527 5807 4561 5835
rect 4589 5807 4623 5835
rect 4651 5807 13437 5835
rect 13465 5807 13499 5835
rect 13527 5807 13561 5835
rect 13589 5807 13623 5835
rect 13651 5807 22437 5835
rect 22465 5807 22499 5835
rect 22527 5807 22561 5835
rect 22589 5807 22623 5835
rect 22651 5807 31437 5835
rect 31465 5807 31499 5835
rect 31527 5807 31561 5835
rect 31589 5807 31623 5835
rect 31651 5807 40437 5835
rect 40465 5807 40499 5835
rect 40527 5807 40561 5835
rect 40589 5807 40623 5835
rect 40651 5807 49437 5835
rect 49465 5807 49499 5835
rect 49527 5807 49561 5835
rect 49589 5807 49623 5835
rect 49651 5807 58437 5835
rect 58465 5807 58499 5835
rect 58527 5807 58561 5835
rect 58589 5807 58623 5835
rect 58651 5807 67437 5835
rect 67465 5807 67499 5835
rect 67527 5807 67561 5835
rect 67589 5807 67623 5835
rect 67651 5807 76437 5835
rect 76465 5807 76499 5835
rect 76527 5807 76561 5835
rect 76589 5807 76623 5835
rect 76651 5807 85437 5835
rect 85465 5807 85499 5835
rect 85527 5807 85561 5835
rect 85589 5807 85623 5835
rect 85651 5807 94437 5835
rect 94465 5807 94499 5835
rect 94527 5807 94561 5835
rect 94589 5807 94623 5835
rect 94651 5807 103437 5835
rect 103465 5807 103499 5835
rect 103527 5807 103561 5835
rect 103589 5807 103623 5835
rect 103651 5807 112437 5835
rect 112465 5807 112499 5835
rect 112527 5807 112561 5835
rect 112589 5807 112623 5835
rect 112651 5807 121437 5835
rect 121465 5807 121499 5835
rect 121527 5807 121561 5835
rect 121589 5807 121623 5835
rect 121651 5807 130437 5835
rect 130465 5807 130499 5835
rect 130527 5807 130561 5835
rect 130589 5807 130623 5835
rect 130651 5807 139437 5835
rect 139465 5807 139499 5835
rect 139527 5807 139561 5835
rect 139589 5807 139623 5835
rect 139651 5807 148437 5835
rect 148465 5807 148499 5835
rect 148527 5807 148561 5835
rect 148589 5807 148623 5835
rect 148651 5807 157437 5835
rect 157465 5807 157499 5835
rect 157527 5807 157561 5835
rect 157589 5807 157623 5835
rect 157651 5807 166437 5835
rect 166465 5807 166499 5835
rect 166527 5807 166561 5835
rect 166589 5807 166623 5835
rect 166651 5807 175437 5835
rect 175465 5807 175499 5835
rect 175527 5807 175561 5835
rect 175589 5807 175623 5835
rect 175651 5807 184437 5835
rect 184465 5807 184499 5835
rect 184527 5807 184561 5835
rect 184589 5807 184623 5835
rect 184651 5807 193437 5835
rect 193465 5807 193499 5835
rect 193527 5807 193561 5835
rect 193589 5807 193623 5835
rect 193651 5807 202437 5835
rect 202465 5807 202499 5835
rect 202527 5807 202561 5835
rect 202589 5807 202623 5835
rect 202651 5807 211437 5835
rect 211465 5807 211499 5835
rect 211527 5807 211561 5835
rect 211589 5807 211623 5835
rect 211651 5807 220437 5835
rect 220465 5807 220499 5835
rect 220527 5807 220561 5835
rect 220589 5807 220623 5835
rect 220651 5807 229437 5835
rect 229465 5807 229499 5835
rect 229527 5807 229561 5835
rect 229589 5807 229623 5835
rect 229651 5807 238437 5835
rect 238465 5807 238499 5835
rect 238527 5807 238561 5835
rect 238589 5807 238623 5835
rect 238651 5807 247437 5835
rect 247465 5807 247499 5835
rect 247527 5807 247561 5835
rect 247589 5807 247623 5835
rect 247651 5807 256437 5835
rect 256465 5807 256499 5835
rect 256527 5807 256561 5835
rect 256589 5807 256623 5835
rect 256651 5807 265437 5835
rect 265465 5807 265499 5835
rect 265527 5807 265561 5835
rect 265589 5807 265623 5835
rect 265651 5807 274437 5835
rect 274465 5807 274499 5835
rect 274527 5807 274561 5835
rect 274589 5807 274623 5835
rect 274651 5807 283437 5835
rect 283465 5807 283499 5835
rect 283527 5807 283561 5835
rect 283589 5807 283623 5835
rect 283651 5807 292437 5835
rect 292465 5807 292499 5835
rect 292527 5807 292561 5835
rect 292589 5807 292623 5835
rect 292651 5807 299736 5835
rect 299764 5807 299798 5835
rect 299826 5807 299860 5835
rect 299888 5807 299922 5835
rect 299950 5807 299998 5835
rect -6 5773 299998 5807
rect -6 5745 42 5773
rect 70 5745 104 5773
rect 132 5745 166 5773
rect 194 5745 228 5773
rect 256 5745 4437 5773
rect 4465 5745 4499 5773
rect 4527 5745 4561 5773
rect 4589 5745 4623 5773
rect 4651 5745 13437 5773
rect 13465 5745 13499 5773
rect 13527 5745 13561 5773
rect 13589 5745 13623 5773
rect 13651 5745 22437 5773
rect 22465 5745 22499 5773
rect 22527 5745 22561 5773
rect 22589 5745 22623 5773
rect 22651 5745 31437 5773
rect 31465 5745 31499 5773
rect 31527 5745 31561 5773
rect 31589 5745 31623 5773
rect 31651 5745 40437 5773
rect 40465 5745 40499 5773
rect 40527 5745 40561 5773
rect 40589 5745 40623 5773
rect 40651 5745 49437 5773
rect 49465 5745 49499 5773
rect 49527 5745 49561 5773
rect 49589 5745 49623 5773
rect 49651 5745 58437 5773
rect 58465 5745 58499 5773
rect 58527 5745 58561 5773
rect 58589 5745 58623 5773
rect 58651 5745 67437 5773
rect 67465 5745 67499 5773
rect 67527 5745 67561 5773
rect 67589 5745 67623 5773
rect 67651 5745 76437 5773
rect 76465 5745 76499 5773
rect 76527 5745 76561 5773
rect 76589 5745 76623 5773
rect 76651 5745 85437 5773
rect 85465 5745 85499 5773
rect 85527 5745 85561 5773
rect 85589 5745 85623 5773
rect 85651 5745 94437 5773
rect 94465 5745 94499 5773
rect 94527 5745 94561 5773
rect 94589 5745 94623 5773
rect 94651 5745 103437 5773
rect 103465 5745 103499 5773
rect 103527 5745 103561 5773
rect 103589 5745 103623 5773
rect 103651 5745 112437 5773
rect 112465 5745 112499 5773
rect 112527 5745 112561 5773
rect 112589 5745 112623 5773
rect 112651 5745 121437 5773
rect 121465 5745 121499 5773
rect 121527 5745 121561 5773
rect 121589 5745 121623 5773
rect 121651 5745 130437 5773
rect 130465 5745 130499 5773
rect 130527 5745 130561 5773
rect 130589 5745 130623 5773
rect 130651 5745 139437 5773
rect 139465 5745 139499 5773
rect 139527 5745 139561 5773
rect 139589 5745 139623 5773
rect 139651 5745 148437 5773
rect 148465 5745 148499 5773
rect 148527 5745 148561 5773
rect 148589 5745 148623 5773
rect 148651 5745 157437 5773
rect 157465 5745 157499 5773
rect 157527 5745 157561 5773
rect 157589 5745 157623 5773
rect 157651 5745 166437 5773
rect 166465 5745 166499 5773
rect 166527 5745 166561 5773
rect 166589 5745 166623 5773
rect 166651 5745 175437 5773
rect 175465 5745 175499 5773
rect 175527 5745 175561 5773
rect 175589 5745 175623 5773
rect 175651 5745 184437 5773
rect 184465 5745 184499 5773
rect 184527 5745 184561 5773
rect 184589 5745 184623 5773
rect 184651 5745 193437 5773
rect 193465 5745 193499 5773
rect 193527 5745 193561 5773
rect 193589 5745 193623 5773
rect 193651 5745 202437 5773
rect 202465 5745 202499 5773
rect 202527 5745 202561 5773
rect 202589 5745 202623 5773
rect 202651 5745 211437 5773
rect 211465 5745 211499 5773
rect 211527 5745 211561 5773
rect 211589 5745 211623 5773
rect 211651 5745 220437 5773
rect 220465 5745 220499 5773
rect 220527 5745 220561 5773
rect 220589 5745 220623 5773
rect 220651 5745 229437 5773
rect 229465 5745 229499 5773
rect 229527 5745 229561 5773
rect 229589 5745 229623 5773
rect 229651 5745 238437 5773
rect 238465 5745 238499 5773
rect 238527 5745 238561 5773
rect 238589 5745 238623 5773
rect 238651 5745 247437 5773
rect 247465 5745 247499 5773
rect 247527 5745 247561 5773
rect 247589 5745 247623 5773
rect 247651 5745 256437 5773
rect 256465 5745 256499 5773
rect 256527 5745 256561 5773
rect 256589 5745 256623 5773
rect 256651 5745 265437 5773
rect 265465 5745 265499 5773
rect 265527 5745 265561 5773
rect 265589 5745 265623 5773
rect 265651 5745 274437 5773
rect 274465 5745 274499 5773
rect 274527 5745 274561 5773
rect 274589 5745 274623 5773
rect 274651 5745 283437 5773
rect 283465 5745 283499 5773
rect 283527 5745 283561 5773
rect 283589 5745 283623 5773
rect 283651 5745 292437 5773
rect 292465 5745 292499 5773
rect 292527 5745 292561 5773
rect 292589 5745 292623 5773
rect 292651 5745 299736 5773
rect 299764 5745 299798 5773
rect 299826 5745 299860 5773
rect 299888 5745 299922 5773
rect 299950 5745 299998 5773
rect -6 5697 299998 5745
rect -6 2959 299998 3007
rect -6 2931 522 2959
rect 550 2931 584 2959
rect 612 2931 646 2959
rect 674 2931 708 2959
rect 736 2931 2577 2959
rect 2605 2931 2639 2959
rect 2667 2931 2701 2959
rect 2729 2931 2763 2959
rect 2791 2931 11577 2959
rect 11605 2931 11639 2959
rect 11667 2931 11701 2959
rect 11729 2931 11763 2959
rect 11791 2931 20577 2959
rect 20605 2931 20639 2959
rect 20667 2931 20701 2959
rect 20729 2931 20763 2959
rect 20791 2931 29577 2959
rect 29605 2931 29639 2959
rect 29667 2931 29701 2959
rect 29729 2931 29763 2959
rect 29791 2931 38577 2959
rect 38605 2931 38639 2959
rect 38667 2931 38701 2959
rect 38729 2931 38763 2959
rect 38791 2931 47577 2959
rect 47605 2931 47639 2959
rect 47667 2931 47701 2959
rect 47729 2931 47763 2959
rect 47791 2931 56577 2959
rect 56605 2931 56639 2959
rect 56667 2931 56701 2959
rect 56729 2931 56763 2959
rect 56791 2931 65577 2959
rect 65605 2931 65639 2959
rect 65667 2931 65701 2959
rect 65729 2931 65763 2959
rect 65791 2931 74577 2959
rect 74605 2931 74639 2959
rect 74667 2931 74701 2959
rect 74729 2931 74763 2959
rect 74791 2931 83577 2959
rect 83605 2931 83639 2959
rect 83667 2931 83701 2959
rect 83729 2931 83763 2959
rect 83791 2931 92577 2959
rect 92605 2931 92639 2959
rect 92667 2931 92701 2959
rect 92729 2931 92763 2959
rect 92791 2931 101577 2959
rect 101605 2931 101639 2959
rect 101667 2931 101701 2959
rect 101729 2931 101763 2959
rect 101791 2931 110577 2959
rect 110605 2931 110639 2959
rect 110667 2931 110701 2959
rect 110729 2931 110763 2959
rect 110791 2931 119577 2959
rect 119605 2931 119639 2959
rect 119667 2931 119701 2959
rect 119729 2931 119763 2959
rect 119791 2931 128577 2959
rect 128605 2931 128639 2959
rect 128667 2931 128701 2959
rect 128729 2931 128763 2959
rect 128791 2931 137577 2959
rect 137605 2931 137639 2959
rect 137667 2931 137701 2959
rect 137729 2931 137763 2959
rect 137791 2931 146577 2959
rect 146605 2931 146639 2959
rect 146667 2931 146701 2959
rect 146729 2931 146763 2959
rect 146791 2931 155577 2959
rect 155605 2931 155639 2959
rect 155667 2931 155701 2959
rect 155729 2931 155763 2959
rect 155791 2931 164577 2959
rect 164605 2931 164639 2959
rect 164667 2931 164701 2959
rect 164729 2931 164763 2959
rect 164791 2931 173577 2959
rect 173605 2931 173639 2959
rect 173667 2931 173701 2959
rect 173729 2931 173763 2959
rect 173791 2931 182577 2959
rect 182605 2931 182639 2959
rect 182667 2931 182701 2959
rect 182729 2931 182763 2959
rect 182791 2931 191577 2959
rect 191605 2931 191639 2959
rect 191667 2931 191701 2959
rect 191729 2931 191763 2959
rect 191791 2931 200577 2959
rect 200605 2931 200639 2959
rect 200667 2931 200701 2959
rect 200729 2931 200763 2959
rect 200791 2931 209577 2959
rect 209605 2931 209639 2959
rect 209667 2931 209701 2959
rect 209729 2931 209763 2959
rect 209791 2931 218577 2959
rect 218605 2931 218639 2959
rect 218667 2931 218701 2959
rect 218729 2931 218763 2959
rect 218791 2931 227577 2959
rect 227605 2931 227639 2959
rect 227667 2931 227701 2959
rect 227729 2931 227763 2959
rect 227791 2931 236577 2959
rect 236605 2931 236639 2959
rect 236667 2931 236701 2959
rect 236729 2931 236763 2959
rect 236791 2931 245577 2959
rect 245605 2931 245639 2959
rect 245667 2931 245701 2959
rect 245729 2931 245763 2959
rect 245791 2931 254577 2959
rect 254605 2931 254639 2959
rect 254667 2931 254701 2959
rect 254729 2931 254763 2959
rect 254791 2931 263577 2959
rect 263605 2931 263639 2959
rect 263667 2931 263701 2959
rect 263729 2931 263763 2959
rect 263791 2931 272577 2959
rect 272605 2931 272639 2959
rect 272667 2931 272701 2959
rect 272729 2931 272763 2959
rect 272791 2931 281577 2959
rect 281605 2931 281639 2959
rect 281667 2931 281701 2959
rect 281729 2931 281763 2959
rect 281791 2931 290577 2959
rect 290605 2931 290639 2959
rect 290667 2931 290701 2959
rect 290729 2931 290763 2959
rect 290791 2931 299256 2959
rect 299284 2931 299318 2959
rect 299346 2931 299380 2959
rect 299408 2931 299442 2959
rect 299470 2931 299998 2959
rect -6 2897 299998 2931
rect -6 2869 522 2897
rect 550 2869 584 2897
rect 612 2869 646 2897
rect 674 2869 708 2897
rect 736 2869 2577 2897
rect 2605 2869 2639 2897
rect 2667 2869 2701 2897
rect 2729 2869 2763 2897
rect 2791 2869 11577 2897
rect 11605 2869 11639 2897
rect 11667 2869 11701 2897
rect 11729 2869 11763 2897
rect 11791 2869 20577 2897
rect 20605 2869 20639 2897
rect 20667 2869 20701 2897
rect 20729 2869 20763 2897
rect 20791 2869 29577 2897
rect 29605 2869 29639 2897
rect 29667 2869 29701 2897
rect 29729 2869 29763 2897
rect 29791 2869 38577 2897
rect 38605 2869 38639 2897
rect 38667 2869 38701 2897
rect 38729 2869 38763 2897
rect 38791 2869 47577 2897
rect 47605 2869 47639 2897
rect 47667 2869 47701 2897
rect 47729 2869 47763 2897
rect 47791 2869 56577 2897
rect 56605 2869 56639 2897
rect 56667 2869 56701 2897
rect 56729 2869 56763 2897
rect 56791 2869 65577 2897
rect 65605 2869 65639 2897
rect 65667 2869 65701 2897
rect 65729 2869 65763 2897
rect 65791 2869 74577 2897
rect 74605 2869 74639 2897
rect 74667 2869 74701 2897
rect 74729 2869 74763 2897
rect 74791 2869 83577 2897
rect 83605 2869 83639 2897
rect 83667 2869 83701 2897
rect 83729 2869 83763 2897
rect 83791 2869 92577 2897
rect 92605 2869 92639 2897
rect 92667 2869 92701 2897
rect 92729 2869 92763 2897
rect 92791 2869 101577 2897
rect 101605 2869 101639 2897
rect 101667 2869 101701 2897
rect 101729 2869 101763 2897
rect 101791 2869 110577 2897
rect 110605 2869 110639 2897
rect 110667 2869 110701 2897
rect 110729 2869 110763 2897
rect 110791 2869 119577 2897
rect 119605 2869 119639 2897
rect 119667 2869 119701 2897
rect 119729 2869 119763 2897
rect 119791 2869 128577 2897
rect 128605 2869 128639 2897
rect 128667 2869 128701 2897
rect 128729 2869 128763 2897
rect 128791 2869 137577 2897
rect 137605 2869 137639 2897
rect 137667 2869 137701 2897
rect 137729 2869 137763 2897
rect 137791 2869 146577 2897
rect 146605 2869 146639 2897
rect 146667 2869 146701 2897
rect 146729 2869 146763 2897
rect 146791 2869 155577 2897
rect 155605 2869 155639 2897
rect 155667 2869 155701 2897
rect 155729 2869 155763 2897
rect 155791 2869 164577 2897
rect 164605 2869 164639 2897
rect 164667 2869 164701 2897
rect 164729 2869 164763 2897
rect 164791 2869 173577 2897
rect 173605 2869 173639 2897
rect 173667 2869 173701 2897
rect 173729 2869 173763 2897
rect 173791 2869 182577 2897
rect 182605 2869 182639 2897
rect 182667 2869 182701 2897
rect 182729 2869 182763 2897
rect 182791 2869 191577 2897
rect 191605 2869 191639 2897
rect 191667 2869 191701 2897
rect 191729 2869 191763 2897
rect 191791 2869 200577 2897
rect 200605 2869 200639 2897
rect 200667 2869 200701 2897
rect 200729 2869 200763 2897
rect 200791 2869 209577 2897
rect 209605 2869 209639 2897
rect 209667 2869 209701 2897
rect 209729 2869 209763 2897
rect 209791 2869 218577 2897
rect 218605 2869 218639 2897
rect 218667 2869 218701 2897
rect 218729 2869 218763 2897
rect 218791 2869 227577 2897
rect 227605 2869 227639 2897
rect 227667 2869 227701 2897
rect 227729 2869 227763 2897
rect 227791 2869 236577 2897
rect 236605 2869 236639 2897
rect 236667 2869 236701 2897
rect 236729 2869 236763 2897
rect 236791 2869 245577 2897
rect 245605 2869 245639 2897
rect 245667 2869 245701 2897
rect 245729 2869 245763 2897
rect 245791 2869 254577 2897
rect 254605 2869 254639 2897
rect 254667 2869 254701 2897
rect 254729 2869 254763 2897
rect 254791 2869 263577 2897
rect 263605 2869 263639 2897
rect 263667 2869 263701 2897
rect 263729 2869 263763 2897
rect 263791 2869 272577 2897
rect 272605 2869 272639 2897
rect 272667 2869 272701 2897
rect 272729 2869 272763 2897
rect 272791 2869 281577 2897
rect 281605 2869 281639 2897
rect 281667 2869 281701 2897
rect 281729 2869 281763 2897
rect 281791 2869 290577 2897
rect 290605 2869 290639 2897
rect 290667 2869 290701 2897
rect 290729 2869 290763 2897
rect 290791 2869 299256 2897
rect 299284 2869 299318 2897
rect 299346 2869 299380 2897
rect 299408 2869 299442 2897
rect 299470 2869 299998 2897
rect -6 2835 299998 2869
rect -6 2807 522 2835
rect 550 2807 584 2835
rect 612 2807 646 2835
rect 674 2807 708 2835
rect 736 2807 2577 2835
rect 2605 2807 2639 2835
rect 2667 2807 2701 2835
rect 2729 2807 2763 2835
rect 2791 2807 11577 2835
rect 11605 2807 11639 2835
rect 11667 2807 11701 2835
rect 11729 2807 11763 2835
rect 11791 2807 20577 2835
rect 20605 2807 20639 2835
rect 20667 2807 20701 2835
rect 20729 2807 20763 2835
rect 20791 2807 29577 2835
rect 29605 2807 29639 2835
rect 29667 2807 29701 2835
rect 29729 2807 29763 2835
rect 29791 2807 38577 2835
rect 38605 2807 38639 2835
rect 38667 2807 38701 2835
rect 38729 2807 38763 2835
rect 38791 2807 47577 2835
rect 47605 2807 47639 2835
rect 47667 2807 47701 2835
rect 47729 2807 47763 2835
rect 47791 2807 56577 2835
rect 56605 2807 56639 2835
rect 56667 2807 56701 2835
rect 56729 2807 56763 2835
rect 56791 2807 65577 2835
rect 65605 2807 65639 2835
rect 65667 2807 65701 2835
rect 65729 2807 65763 2835
rect 65791 2807 74577 2835
rect 74605 2807 74639 2835
rect 74667 2807 74701 2835
rect 74729 2807 74763 2835
rect 74791 2807 83577 2835
rect 83605 2807 83639 2835
rect 83667 2807 83701 2835
rect 83729 2807 83763 2835
rect 83791 2807 92577 2835
rect 92605 2807 92639 2835
rect 92667 2807 92701 2835
rect 92729 2807 92763 2835
rect 92791 2807 101577 2835
rect 101605 2807 101639 2835
rect 101667 2807 101701 2835
rect 101729 2807 101763 2835
rect 101791 2807 110577 2835
rect 110605 2807 110639 2835
rect 110667 2807 110701 2835
rect 110729 2807 110763 2835
rect 110791 2807 119577 2835
rect 119605 2807 119639 2835
rect 119667 2807 119701 2835
rect 119729 2807 119763 2835
rect 119791 2807 128577 2835
rect 128605 2807 128639 2835
rect 128667 2807 128701 2835
rect 128729 2807 128763 2835
rect 128791 2807 137577 2835
rect 137605 2807 137639 2835
rect 137667 2807 137701 2835
rect 137729 2807 137763 2835
rect 137791 2807 146577 2835
rect 146605 2807 146639 2835
rect 146667 2807 146701 2835
rect 146729 2807 146763 2835
rect 146791 2807 155577 2835
rect 155605 2807 155639 2835
rect 155667 2807 155701 2835
rect 155729 2807 155763 2835
rect 155791 2807 164577 2835
rect 164605 2807 164639 2835
rect 164667 2807 164701 2835
rect 164729 2807 164763 2835
rect 164791 2807 173577 2835
rect 173605 2807 173639 2835
rect 173667 2807 173701 2835
rect 173729 2807 173763 2835
rect 173791 2807 182577 2835
rect 182605 2807 182639 2835
rect 182667 2807 182701 2835
rect 182729 2807 182763 2835
rect 182791 2807 191577 2835
rect 191605 2807 191639 2835
rect 191667 2807 191701 2835
rect 191729 2807 191763 2835
rect 191791 2807 200577 2835
rect 200605 2807 200639 2835
rect 200667 2807 200701 2835
rect 200729 2807 200763 2835
rect 200791 2807 209577 2835
rect 209605 2807 209639 2835
rect 209667 2807 209701 2835
rect 209729 2807 209763 2835
rect 209791 2807 218577 2835
rect 218605 2807 218639 2835
rect 218667 2807 218701 2835
rect 218729 2807 218763 2835
rect 218791 2807 227577 2835
rect 227605 2807 227639 2835
rect 227667 2807 227701 2835
rect 227729 2807 227763 2835
rect 227791 2807 236577 2835
rect 236605 2807 236639 2835
rect 236667 2807 236701 2835
rect 236729 2807 236763 2835
rect 236791 2807 245577 2835
rect 245605 2807 245639 2835
rect 245667 2807 245701 2835
rect 245729 2807 245763 2835
rect 245791 2807 254577 2835
rect 254605 2807 254639 2835
rect 254667 2807 254701 2835
rect 254729 2807 254763 2835
rect 254791 2807 263577 2835
rect 263605 2807 263639 2835
rect 263667 2807 263701 2835
rect 263729 2807 263763 2835
rect 263791 2807 272577 2835
rect 272605 2807 272639 2835
rect 272667 2807 272701 2835
rect 272729 2807 272763 2835
rect 272791 2807 281577 2835
rect 281605 2807 281639 2835
rect 281667 2807 281701 2835
rect 281729 2807 281763 2835
rect 281791 2807 290577 2835
rect 290605 2807 290639 2835
rect 290667 2807 290701 2835
rect 290729 2807 290763 2835
rect 290791 2807 299256 2835
rect 299284 2807 299318 2835
rect 299346 2807 299380 2835
rect 299408 2807 299442 2835
rect 299470 2807 299998 2835
rect -6 2773 299998 2807
rect -6 2745 522 2773
rect 550 2745 584 2773
rect 612 2745 646 2773
rect 674 2745 708 2773
rect 736 2745 2577 2773
rect 2605 2745 2639 2773
rect 2667 2745 2701 2773
rect 2729 2745 2763 2773
rect 2791 2745 11577 2773
rect 11605 2745 11639 2773
rect 11667 2745 11701 2773
rect 11729 2745 11763 2773
rect 11791 2745 20577 2773
rect 20605 2745 20639 2773
rect 20667 2745 20701 2773
rect 20729 2745 20763 2773
rect 20791 2745 29577 2773
rect 29605 2745 29639 2773
rect 29667 2745 29701 2773
rect 29729 2745 29763 2773
rect 29791 2745 38577 2773
rect 38605 2745 38639 2773
rect 38667 2745 38701 2773
rect 38729 2745 38763 2773
rect 38791 2745 47577 2773
rect 47605 2745 47639 2773
rect 47667 2745 47701 2773
rect 47729 2745 47763 2773
rect 47791 2745 56577 2773
rect 56605 2745 56639 2773
rect 56667 2745 56701 2773
rect 56729 2745 56763 2773
rect 56791 2745 65577 2773
rect 65605 2745 65639 2773
rect 65667 2745 65701 2773
rect 65729 2745 65763 2773
rect 65791 2745 74577 2773
rect 74605 2745 74639 2773
rect 74667 2745 74701 2773
rect 74729 2745 74763 2773
rect 74791 2745 83577 2773
rect 83605 2745 83639 2773
rect 83667 2745 83701 2773
rect 83729 2745 83763 2773
rect 83791 2745 92577 2773
rect 92605 2745 92639 2773
rect 92667 2745 92701 2773
rect 92729 2745 92763 2773
rect 92791 2745 101577 2773
rect 101605 2745 101639 2773
rect 101667 2745 101701 2773
rect 101729 2745 101763 2773
rect 101791 2745 110577 2773
rect 110605 2745 110639 2773
rect 110667 2745 110701 2773
rect 110729 2745 110763 2773
rect 110791 2745 119577 2773
rect 119605 2745 119639 2773
rect 119667 2745 119701 2773
rect 119729 2745 119763 2773
rect 119791 2745 128577 2773
rect 128605 2745 128639 2773
rect 128667 2745 128701 2773
rect 128729 2745 128763 2773
rect 128791 2745 137577 2773
rect 137605 2745 137639 2773
rect 137667 2745 137701 2773
rect 137729 2745 137763 2773
rect 137791 2745 146577 2773
rect 146605 2745 146639 2773
rect 146667 2745 146701 2773
rect 146729 2745 146763 2773
rect 146791 2745 155577 2773
rect 155605 2745 155639 2773
rect 155667 2745 155701 2773
rect 155729 2745 155763 2773
rect 155791 2745 164577 2773
rect 164605 2745 164639 2773
rect 164667 2745 164701 2773
rect 164729 2745 164763 2773
rect 164791 2745 173577 2773
rect 173605 2745 173639 2773
rect 173667 2745 173701 2773
rect 173729 2745 173763 2773
rect 173791 2745 182577 2773
rect 182605 2745 182639 2773
rect 182667 2745 182701 2773
rect 182729 2745 182763 2773
rect 182791 2745 191577 2773
rect 191605 2745 191639 2773
rect 191667 2745 191701 2773
rect 191729 2745 191763 2773
rect 191791 2745 200577 2773
rect 200605 2745 200639 2773
rect 200667 2745 200701 2773
rect 200729 2745 200763 2773
rect 200791 2745 209577 2773
rect 209605 2745 209639 2773
rect 209667 2745 209701 2773
rect 209729 2745 209763 2773
rect 209791 2745 218577 2773
rect 218605 2745 218639 2773
rect 218667 2745 218701 2773
rect 218729 2745 218763 2773
rect 218791 2745 227577 2773
rect 227605 2745 227639 2773
rect 227667 2745 227701 2773
rect 227729 2745 227763 2773
rect 227791 2745 236577 2773
rect 236605 2745 236639 2773
rect 236667 2745 236701 2773
rect 236729 2745 236763 2773
rect 236791 2745 245577 2773
rect 245605 2745 245639 2773
rect 245667 2745 245701 2773
rect 245729 2745 245763 2773
rect 245791 2745 254577 2773
rect 254605 2745 254639 2773
rect 254667 2745 254701 2773
rect 254729 2745 254763 2773
rect 254791 2745 263577 2773
rect 263605 2745 263639 2773
rect 263667 2745 263701 2773
rect 263729 2745 263763 2773
rect 263791 2745 272577 2773
rect 272605 2745 272639 2773
rect 272667 2745 272701 2773
rect 272729 2745 272763 2773
rect 272791 2745 281577 2773
rect 281605 2745 281639 2773
rect 281667 2745 281701 2773
rect 281729 2745 281763 2773
rect 281791 2745 290577 2773
rect 290605 2745 290639 2773
rect 290667 2745 290701 2773
rect 290729 2745 290763 2773
rect 290791 2745 299256 2773
rect 299284 2745 299318 2773
rect 299346 2745 299380 2773
rect 299408 2745 299442 2773
rect 299470 2745 299998 2773
rect -6 2697 299998 2745
rect 474 904 299518 952
rect 474 876 522 904
rect 550 876 584 904
rect 612 876 646 904
rect 674 876 708 904
rect 736 876 2577 904
rect 2605 876 2639 904
rect 2667 876 2701 904
rect 2729 876 2763 904
rect 2791 876 11577 904
rect 11605 876 11639 904
rect 11667 876 11701 904
rect 11729 876 11763 904
rect 11791 876 20577 904
rect 20605 876 20639 904
rect 20667 876 20701 904
rect 20729 876 20763 904
rect 20791 876 29577 904
rect 29605 876 29639 904
rect 29667 876 29701 904
rect 29729 876 29763 904
rect 29791 876 38577 904
rect 38605 876 38639 904
rect 38667 876 38701 904
rect 38729 876 38763 904
rect 38791 876 47577 904
rect 47605 876 47639 904
rect 47667 876 47701 904
rect 47729 876 47763 904
rect 47791 876 56577 904
rect 56605 876 56639 904
rect 56667 876 56701 904
rect 56729 876 56763 904
rect 56791 876 65577 904
rect 65605 876 65639 904
rect 65667 876 65701 904
rect 65729 876 65763 904
rect 65791 876 74577 904
rect 74605 876 74639 904
rect 74667 876 74701 904
rect 74729 876 74763 904
rect 74791 876 83577 904
rect 83605 876 83639 904
rect 83667 876 83701 904
rect 83729 876 83763 904
rect 83791 876 92577 904
rect 92605 876 92639 904
rect 92667 876 92701 904
rect 92729 876 92763 904
rect 92791 876 101577 904
rect 101605 876 101639 904
rect 101667 876 101701 904
rect 101729 876 101763 904
rect 101791 876 110577 904
rect 110605 876 110639 904
rect 110667 876 110701 904
rect 110729 876 110763 904
rect 110791 876 119577 904
rect 119605 876 119639 904
rect 119667 876 119701 904
rect 119729 876 119763 904
rect 119791 876 128577 904
rect 128605 876 128639 904
rect 128667 876 128701 904
rect 128729 876 128763 904
rect 128791 876 137577 904
rect 137605 876 137639 904
rect 137667 876 137701 904
rect 137729 876 137763 904
rect 137791 876 146577 904
rect 146605 876 146639 904
rect 146667 876 146701 904
rect 146729 876 146763 904
rect 146791 876 155577 904
rect 155605 876 155639 904
rect 155667 876 155701 904
rect 155729 876 155763 904
rect 155791 876 164577 904
rect 164605 876 164639 904
rect 164667 876 164701 904
rect 164729 876 164763 904
rect 164791 876 173577 904
rect 173605 876 173639 904
rect 173667 876 173701 904
rect 173729 876 173763 904
rect 173791 876 182577 904
rect 182605 876 182639 904
rect 182667 876 182701 904
rect 182729 876 182763 904
rect 182791 876 191577 904
rect 191605 876 191639 904
rect 191667 876 191701 904
rect 191729 876 191763 904
rect 191791 876 200577 904
rect 200605 876 200639 904
rect 200667 876 200701 904
rect 200729 876 200763 904
rect 200791 876 209577 904
rect 209605 876 209639 904
rect 209667 876 209701 904
rect 209729 876 209763 904
rect 209791 876 218577 904
rect 218605 876 218639 904
rect 218667 876 218701 904
rect 218729 876 218763 904
rect 218791 876 227577 904
rect 227605 876 227639 904
rect 227667 876 227701 904
rect 227729 876 227763 904
rect 227791 876 236577 904
rect 236605 876 236639 904
rect 236667 876 236701 904
rect 236729 876 236763 904
rect 236791 876 245577 904
rect 245605 876 245639 904
rect 245667 876 245701 904
rect 245729 876 245763 904
rect 245791 876 254577 904
rect 254605 876 254639 904
rect 254667 876 254701 904
rect 254729 876 254763 904
rect 254791 876 263577 904
rect 263605 876 263639 904
rect 263667 876 263701 904
rect 263729 876 263763 904
rect 263791 876 272577 904
rect 272605 876 272639 904
rect 272667 876 272701 904
rect 272729 876 272763 904
rect 272791 876 281577 904
rect 281605 876 281639 904
rect 281667 876 281701 904
rect 281729 876 281763 904
rect 281791 876 290577 904
rect 290605 876 290639 904
rect 290667 876 290701 904
rect 290729 876 290763 904
rect 290791 876 299256 904
rect 299284 876 299318 904
rect 299346 876 299380 904
rect 299408 876 299442 904
rect 299470 876 299518 904
rect 474 842 299518 876
rect 474 814 522 842
rect 550 814 584 842
rect 612 814 646 842
rect 674 814 708 842
rect 736 814 2577 842
rect 2605 814 2639 842
rect 2667 814 2701 842
rect 2729 814 2763 842
rect 2791 814 11577 842
rect 11605 814 11639 842
rect 11667 814 11701 842
rect 11729 814 11763 842
rect 11791 814 20577 842
rect 20605 814 20639 842
rect 20667 814 20701 842
rect 20729 814 20763 842
rect 20791 814 29577 842
rect 29605 814 29639 842
rect 29667 814 29701 842
rect 29729 814 29763 842
rect 29791 814 38577 842
rect 38605 814 38639 842
rect 38667 814 38701 842
rect 38729 814 38763 842
rect 38791 814 47577 842
rect 47605 814 47639 842
rect 47667 814 47701 842
rect 47729 814 47763 842
rect 47791 814 56577 842
rect 56605 814 56639 842
rect 56667 814 56701 842
rect 56729 814 56763 842
rect 56791 814 65577 842
rect 65605 814 65639 842
rect 65667 814 65701 842
rect 65729 814 65763 842
rect 65791 814 74577 842
rect 74605 814 74639 842
rect 74667 814 74701 842
rect 74729 814 74763 842
rect 74791 814 83577 842
rect 83605 814 83639 842
rect 83667 814 83701 842
rect 83729 814 83763 842
rect 83791 814 92577 842
rect 92605 814 92639 842
rect 92667 814 92701 842
rect 92729 814 92763 842
rect 92791 814 101577 842
rect 101605 814 101639 842
rect 101667 814 101701 842
rect 101729 814 101763 842
rect 101791 814 110577 842
rect 110605 814 110639 842
rect 110667 814 110701 842
rect 110729 814 110763 842
rect 110791 814 119577 842
rect 119605 814 119639 842
rect 119667 814 119701 842
rect 119729 814 119763 842
rect 119791 814 128577 842
rect 128605 814 128639 842
rect 128667 814 128701 842
rect 128729 814 128763 842
rect 128791 814 137577 842
rect 137605 814 137639 842
rect 137667 814 137701 842
rect 137729 814 137763 842
rect 137791 814 146577 842
rect 146605 814 146639 842
rect 146667 814 146701 842
rect 146729 814 146763 842
rect 146791 814 155577 842
rect 155605 814 155639 842
rect 155667 814 155701 842
rect 155729 814 155763 842
rect 155791 814 164577 842
rect 164605 814 164639 842
rect 164667 814 164701 842
rect 164729 814 164763 842
rect 164791 814 173577 842
rect 173605 814 173639 842
rect 173667 814 173701 842
rect 173729 814 173763 842
rect 173791 814 182577 842
rect 182605 814 182639 842
rect 182667 814 182701 842
rect 182729 814 182763 842
rect 182791 814 191577 842
rect 191605 814 191639 842
rect 191667 814 191701 842
rect 191729 814 191763 842
rect 191791 814 200577 842
rect 200605 814 200639 842
rect 200667 814 200701 842
rect 200729 814 200763 842
rect 200791 814 209577 842
rect 209605 814 209639 842
rect 209667 814 209701 842
rect 209729 814 209763 842
rect 209791 814 218577 842
rect 218605 814 218639 842
rect 218667 814 218701 842
rect 218729 814 218763 842
rect 218791 814 227577 842
rect 227605 814 227639 842
rect 227667 814 227701 842
rect 227729 814 227763 842
rect 227791 814 236577 842
rect 236605 814 236639 842
rect 236667 814 236701 842
rect 236729 814 236763 842
rect 236791 814 245577 842
rect 245605 814 245639 842
rect 245667 814 245701 842
rect 245729 814 245763 842
rect 245791 814 254577 842
rect 254605 814 254639 842
rect 254667 814 254701 842
rect 254729 814 254763 842
rect 254791 814 263577 842
rect 263605 814 263639 842
rect 263667 814 263701 842
rect 263729 814 263763 842
rect 263791 814 272577 842
rect 272605 814 272639 842
rect 272667 814 272701 842
rect 272729 814 272763 842
rect 272791 814 281577 842
rect 281605 814 281639 842
rect 281667 814 281701 842
rect 281729 814 281763 842
rect 281791 814 290577 842
rect 290605 814 290639 842
rect 290667 814 290701 842
rect 290729 814 290763 842
rect 290791 814 299256 842
rect 299284 814 299318 842
rect 299346 814 299380 842
rect 299408 814 299442 842
rect 299470 814 299518 842
rect 474 780 299518 814
rect 474 752 522 780
rect 550 752 584 780
rect 612 752 646 780
rect 674 752 708 780
rect 736 752 2577 780
rect 2605 752 2639 780
rect 2667 752 2701 780
rect 2729 752 2763 780
rect 2791 752 11577 780
rect 11605 752 11639 780
rect 11667 752 11701 780
rect 11729 752 11763 780
rect 11791 752 20577 780
rect 20605 752 20639 780
rect 20667 752 20701 780
rect 20729 752 20763 780
rect 20791 752 29577 780
rect 29605 752 29639 780
rect 29667 752 29701 780
rect 29729 752 29763 780
rect 29791 752 38577 780
rect 38605 752 38639 780
rect 38667 752 38701 780
rect 38729 752 38763 780
rect 38791 752 47577 780
rect 47605 752 47639 780
rect 47667 752 47701 780
rect 47729 752 47763 780
rect 47791 752 56577 780
rect 56605 752 56639 780
rect 56667 752 56701 780
rect 56729 752 56763 780
rect 56791 752 65577 780
rect 65605 752 65639 780
rect 65667 752 65701 780
rect 65729 752 65763 780
rect 65791 752 74577 780
rect 74605 752 74639 780
rect 74667 752 74701 780
rect 74729 752 74763 780
rect 74791 752 83577 780
rect 83605 752 83639 780
rect 83667 752 83701 780
rect 83729 752 83763 780
rect 83791 752 92577 780
rect 92605 752 92639 780
rect 92667 752 92701 780
rect 92729 752 92763 780
rect 92791 752 101577 780
rect 101605 752 101639 780
rect 101667 752 101701 780
rect 101729 752 101763 780
rect 101791 752 110577 780
rect 110605 752 110639 780
rect 110667 752 110701 780
rect 110729 752 110763 780
rect 110791 752 119577 780
rect 119605 752 119639 780
rect 119667 752 119701 780
rect 119729 752 119763 780
rect 119791 752 128577 780
rect 128605 752 128639 780
rect 128667 752 128701 780
rect 128729 752 128763 780
rect 128791 752 137577 780
rect 137605 752 137639 780
rect 137667 752 137701 780
rect 137729 752 137763 780
rect 137791 752 146577 780
rect 146605 752 146639 780
rect 146667 752 146701 780
rect 146729 752 146763 780
rect 146791 752 155577 780
rect 155605 752 155639 780
rect 155667 752 155701 780
rect 155729 752 155763 780
rect 155791 752 164577 780
rect 164605 752 164639 780
rect 164667 752 164701 780
rect 164729 752 164763 780
rect 164791 752 173577 780
rect 173605 752 173639 780
rect 173667 752 173701 780
rect 173729 752 173763 780
rect 173791 752 182577 780
rect 182605 752 182639 780
rect 182667 752 182701 780
rect 182729 752 182763 780
rect 182791 752 191577 780
rect 191605 752 191639 780
rect 191667 752 191701 780
rect 191729 752 191763 780
rect 191791 752 200577 780
rect 200605 752 200639 780
rect 200667 752 200701 780
rect 200729 752 200763 780
rect 200791 752 209577 780
rect 209605 752 209639 780
rect 209667 752 209701 780
rect 209729 752 209763 780
rect 209791 752 218577 780
rect 218605 752 218639 780
rect 218667 752 218701 780
rect 218729 752 218763 780
rect 218791 752 227577 780
rect 227605 752 227639 780
rect 227667 752 227701 780
rect 227729 752 227763 780
rect 227791 752 236577 780
rect 236605 752 236639 780
rect 236667 752 236701 780
rect 236729 752 236763 780
rect 236791 752 245577 780
rect 245605 752 245639 780
rect 245667 752 245701 780
rect 245729 752 245763 780
rect 245791 752 254577 780
rect 254605 752 254639 780
rect 254667 752 254701 780
rect 254729 752 254763 780
rect 254791 752 263577 780
rect 263605 752 263639 780
rect 263667 752 263701 780
rect 263729 752 263763 780
rect 263791 752 272577 780
rect 272605 752 272639 780
rect 272667 752 272701 780
rect 272729 752 272763 780
rect 272791 752 281577 780
rect 281605 752 281639 780
rect 281667 752 281701 780
rect 281729 752 281763 780
rect 281791 752 290577 780
rect 290605 752 290639 780
rect 290667 752 290701 780
rect 290729 752 290763 780
rect 290791 752 299256 780
rect 299284 752 299318 780
rect 299346 752 299380 780
rect 299408 752 299442 780
rect 299470 752 299518 780
rect 474 718 299518 752
rect 474 690 522 718
rect 550 690 584 718
rect 612 690 646 718
rect 674 690 708 718
rect 736 690 2577 718
rect 2605 690 2639 718
rect 2667 690 2701 718
rect 2729 690 2763 718
rect 2791 690 11577 718
rect 11605 690 11639 718
rect 11667 690 11701 718
rect 11729 690 11763 718
rect 11791 690 20577 718
rect 20605 690 20639 718
rect 20667 690 20701 718
rect 20729 690 20763 718
rect 20791 690 29577 718
rect 29605 690 29639 718
rect 29667 690 29701 718
rect 29729 690 29763 718
rect 29791 690 38577 718
rect 38605 690 38639 718
rect 38667 690 38701 718
rect 38729 690 38763 718
rect 38791 690 47577 718
rect 47605 690 47639 718
rect 47667 690 47701 718
rect 47729 690 47763 718
rect 47791 690 56577 718
rect 56605 690 56639 718
rect 56667 690 56701 718
rect 56729 690 56763 718
rect 56791 690 65577 718
rect 65605 690 65639 718
rect 65667 690 65701 718
rect 65729 690 65763 718
rect 65791 690 74577 718
rect 74605 690 74639 718
rect 74667 690 74701 718
rect 74729 690 74763 718
rect 74791 690 83577 718
rect 83605 690 83639 718
rect 83667 690 83701 718
rect 83729 690 83763 718
rect 83791 690 92577 718
rect 92605 690 92639 718
rect 92667 690 92701 718
rect 92729 690 92763 718
rect 92791 690 101577 718
rect 101605 690 101639 718
rect 101667 690 101701 718
rect 101729 690 101763 718
rect 101791 690 110577 718
rect 110605 690 110639 718
rect 110667 690 110701 718
rect 110729 690 110763 718
rect 110791 690 119577 718
rect 119605 690 119639 718
rect 119667 690 119701 718
rect 119729 690 119763 718
rect 119791 690 128577 718
rect 128605 690 128639 718
rect 128667 690 128701 718
rect 128729 690 128763 718
rect 128791 690 137577 718
rect 137605 690 137639 718
rect 137667 690 137701 718
rect 137729 690 137763 718
rect 137791 690 146577 718
rect 146605 690 146639 718
rect 146667 690 146701 718
rect 146729 690 146763 718
rect 146791 690 155577 718
rect 155605 690 155639 718
rect 155667 690 155701 718
rect 155729 690 155763 718
rect 155791 690 164577 718
rect 164605 690 164639 718
rect 164667 690 164701 718
rect 164729 690 164763 718
rect 164791 690 173577 718
rect 173605 690 173639 718
rect 173667 690 173701 718
rect 173729 690 173763 718
rect 173791 690 182577 718
rect 182605 690 182639 718
rect 182667 690 182701 718
rect 182729 690 182763 718
rect 182791 690 191577 718
rect 191605 690 191639 718
rect 191667 690 191701 718
rect 191729 690 191763 718
rect 191791 690 200577 718
rect 200605 690 200639 718
rect 200667 690 200701 718
rect 200729 690 200763 718
rect 200791 690 209577 718
rect 209605 690 209639 718
rect 209667 690 209701 718
rect 209729 690 209763 718
rect 209791 690 218577 718
rect 218605 690 218639 718
rect 218667 690 218701 718
rect 218729 690 218763 718
rect 218791 690 227577 718
rect 227605 690 227639 718
rect 227667 690 227701 718
rect 227729 690 227763 718
rect 227791 690 236577 718
rect 236605 690 236639 718
rect 236667 690 236701 718
rect 236729 690 236763 718
rect 236791 690 245577 718
rect 245605 690 245639 718
rect 245667 690 245701 718
rect 245729 690 245763 718
rect 245791 690 254577 718
rect 254605 690 254639 718
rect 254667 690 254701 718
rect 254729 690 254763 718
rect 254791 690 263577 718
rect 263605 690 263639 718
rect 263667 690 263701 718
rect 263729 690 263763 718
rect 263791 690 272577 718
rect 272605 690 272639 718
rect 272667 690 272701 718
rect 272729 690 272763 718
rect 272791 690 281577 718
rect 281605 690 281639 718
rect 281667 690 281701 718
rect 281729 690 281763 718
rect 281791 690 290577 718
rect 290605 690 290639 718
rect 290667 690 290701 718
rect 290729 690 290763 718
rect 290791 690 299256 718
rect 299284 690 299318 718
rect 299346 690 299380 718
rect 299408 690 299442 718
rect 299470 690 299518 718
rect 474 642 299518 690
rect -6 424 299998 472
rect -6 396 42 424
rect 70 396 104 424
rect 132 396 166 424
rect 194 396 228 424
rect 256 396 4437 424
rect 4465 396 4499 424
rect 4527 396 4561 424
rect 4589 396 4623 424
rect 4651 396 13437 424
rect 13465 396 13499 424
rect 13527 396 13561 424
rect 13589 396 13623 424
rect 13651 396 22437 424
rect 22465 396 22499 424
rect 22527 396 22561 424
rect 22589 396 22623 424
rect 22651 396 31437 424
rect 31465 396 31499 424
rect 31527 396 31561 424
rect 31589 396 31623 424
rect 31651 396 40437 424
rect 40465 396 40499 424
rect 40527 396 40561 424
rect 40589 396 40623 424
rect 40651 396 49437 424
rect 49465 396 49499 424
rect 49527 396 49561 424
rect 49589 396 49623 424
rect 49651 396 58437 424
rect 58465 396 58499 424
rect 58527 396 58561 424
rect 58589 396 58623 424
rect 58651 396 67437 424
rect 67465 396 67499 424
rect 67527 396 67561 424
rect 67589 396 67623 424
rect 67651 396 76437 424
rect 76465 396 76499 424
rect 76527 396 76561 424
rect 76589 396 76623 424
rect 76651 396 85437 424
rect 85465 396 85499 424
rect 85527 396 85561 424
rect 85589 396 85623 424
rect 85651 396 94437 424
rect 94465 396 94499 424
rect 94527 396 94561 424
rect 94589 396 94623 424
rect 94651 396 103437 424
rect 103465 396 103499 424
rect 103527 396 103561 424
rect 103589 396 103623 424
rect 103651 396 112437 424
rect 112465 396 112499 424
rect 112527 396 112561 424
rect 112589 396 112623 424
rect 112651 396 121437 424
rect 121465 396 121499 424
rect 121527 396 121561 424
rect 121589 396 121623 424
rect 121651 396 130437 424
rect 130465 396 130499 424
rect 130527 396 130561 424
rect 130589 396 130623 424
rect 130651 396 139437 424
rect 139465 396 139499 424
rect 139527 396 139561 424
rect 139589 396 139623 424
rect 139651 396 148437 424
rect 148465 396 148499 424
rect 148527 396 148561 424
rect 148589 396 148623 424
rect 148651 396 157437 424
rect 157465 396 157499 424
rect 157527 396 157561 424
rect 157589 396 157623 424
rect 157651 396 166437 424
rect 166465 396 166499 424
rect 166527 396 166561 424
rect 166589 396 166623 424
rect 166651 396 175437 424
rect 175465 396 175499 424
rect 175527 396 175561 424
rect 175589 396 175623 424
rect 175651 396 184437 424
rect 184465 396 184499 424
rect 184527 396 184561 424
rect 184589 396 184623 424
rect 184651 396 193437 424
rect 193465 396 193499 424
rect 193527 396 193561 424
rect 193589 396 193623 424
rect 193651 396 202437 424
rect 202465 396 202499 424
rect 202527 396 202561 424
rect 202589 396 202623 424
rect 202651 396 211437 424
rect 211465 396 211499 424
rect 211527 396 211561 424
rect 211589 396 211623 424
rect 211651 396 220437 424
rect 220465 396 220499 424
rect 220527 396 220561 424
rect 220589 396 220623 424
rect 220651 396 229437 424
rect 229465 396 229499 424
rect 229527 396 229561 424
rect 229589 396 229623 424
rect 229651 396 238437 424
rect 238465 396 238499 424
rect 238527 396 238561 424
rect 238589 396 238623 424
rect 238651 396 247437 424
rect 247465 396 247499 424
rect 247527 396 247561 424
rect 247589 396 247623 424
rect 247651 396 256437 424
rect 256465 396 256499 424
rect 256527 396 256561 424
rect 256589 396 256623 424
rect 256651 396 265437 424
rect 265465 396 265499 424
rect 265527 396 265561 424
rect 265589 396 265623 424
rect 265651 396 274437 424
rect 274465 396 274499 424
rect 274527 396 274561 424
rect 274589 396 274623 424
rect 274651 396 283437 424
rect 283465 396 283499 424
rect 283527 396 283561 424
rect 283589 396 283623 424
rect 283651 396 292437 424
rect 292465 396 292499 424
rect 292527 396 292561 424
rect 292589 396 292623 424
rect 292651 396 299736 424
rect 299764 396 299798 424
rect 299826 396 299860 424
rect 299888 396 299922 424
rect 299950 396 299998 424
rect -6 362 299998 396
rect -6 334 42 362
rect 70 334 104 362
rect 132 334 166 362
rect 194 334 228 362
rect 256 334 4437 362
rect 4465 334 4499 362
rect 4527 334 4561 362
rect 4589 334 4623 362
rect 4651 334 13437 362
rect 13465 334 13499 362
rect 13527 334 13561 362
rect 13589 334 13623 362
rect 13651 334 22437 362
rect 22465 334 22499 362
rect 22527 334 22561 362
rect 22589 334 22623 362
rect 22651 334 31437 362
rect 31465 334 31499 362
rect 31527 334 31561 362
rect 31589 334 31623 362
rect 31651 334 40437 362
rect 40465 334 40499 362
rect 40527 334 40561 362
rect 40589 334 40623 362
rect 40651 334 49437 362
rect 49465 334 49499 362
rect 49527 334 49561 362
rect 49589 334 49623 362
rect 49651 334 58437 362
rect 58465 334 58499 362
rect 58527 334 58561 362
rect 58589 334 58623 362
rect 58651 334 67437 362
rect 67465 334 67499 362
rect 67527 334 67561 362
rect 67589 334 67623 362
rect 67651 334 76437 362
rect 76465 334 76499 362
rect 76527 334 76561 362
rect 76589 334 76623 362
rect 76651 334 85437 362
rect 85465 334 85499 362
rect 85527 334 85561 362
rect 85589 334 85623 362
rect 85651 334 94437 362
rect 94465 334 94499 362
rect 94527 334 94561 362
rect 94589 334 94623 362
rect 94651 334 103437 362
rect 103465 334 103499 362
rect 103527 334 103561 362
rect 103589 334 103623 362
rect 103651 334 112437 362
rect 112465 334 112499 362
rect 112527 334 112561 362
rect 112589 334 112623 362
rect 112651 334 121437 362
rect 121465 334 121499 362
rect 121527 334 121561 362
rect 121589 334 121623 362
rect 121651 334 130437 362
rect 130465 334 130499 362
rect 130527 334 130561 362
rect 130589 334 130623 362
rect 130651 334 139437 362
rect 139465 334 139499 362
rect 139527 334 139561 362
rect 139589 334 139623 362
rect 139651 334 148437 362
rect 148465 334 148499 362
rect 148527 334 148561 362
rect 148589 334 148623 362
rect 148651 334 157437 362
rect 157465 334 157499 362
rect 157527 334 157561 362
rect 157589 334 157623 362
rect 157651 334 166437 362
rect 166465 334 166499 362
rect 166527 334 166561 362
rect 166589 334 166623 362
rect 166651 334 175437 362
rect 175465 334 175499 362
rect 175527 334 175561 362
rect 175589 334 175623 362
rect 175651 334 184437 362
rect 184465 334 184499 362
rect 184527 334 184561 362
rect 184589 334 184623 362
rect 184651 334 193437 362
rect 193465 334 193499 362
rect 193527 334 193561 362
rect 193589 334 193623 362
rect 193651 334 202437 362
rect 202465 334 202499 362
rect 202527 334 202561 362
rect 202589 334 202623 362
rect 202651 334 211437 362
rect 211465 334 211499 362
rect 211527 334 211561 362
rect 211589 334 211623 362
rect 211651 334 220437 362
rect 220465 334 220499 362
rect 220527 334 220561 362
rect 220589 334 220623 362
rect 220651 334 229437 362
rect 229465 334 229499 362
rect 229527 334 229561 362
rect 229589 334 229623 362
rect 229651 334 238437 362
rect 238465 334 238499 362
rect 238527 334 238561 362
rect 238589 334 238623 362
rect 238651 334 247437 362
rect 247465 334 247499 362
rect 247527 334 247561 362
rect 247589 334 247623 362
rect 247651 334 256437 362
rect 256465 334 256499 362
rect 256527 334 256561 362
rect 256589 334 256623 362
rect 256651 334 265437 362
rect 265465 334 265499 362
rect 265527 334 265561 362
rect 265589 334 265623 362
rect 265651 334 274437 362
rect 274465 334 274499 362
rect 274527 334 274561 362
rect 274589 334 274623 362
rect 274651 334 283437 362
rect 283465 334 283499 362
rect 283527 334 283561 362
rect 283589 334 283623 362
rect 283651 334 292437 362
rect 292465 334 292499 362
rect 292527 334 292561 362
rect 292589 334 292623 362
rect 292651 334 299736 362
rect 299764 334 299798 362
rect 299826 334 299860 362
rect 299888 334 299922 362
rect 299950 334 299998 362
rect -6 300 299998 334
rect -6 272 42 300
rect 70 272 104 300
rect 132 272 166 300
rect 194 272 228 300
rect 256 272 4437 300
rect 4465 272 4499 300
rect 4527 272 4561 300
rect 4589 272 4623 300
rect 4651 272 13437 300
rect 13465 272 13499 300
rect 13527 272 13561 300
rect 13589 272 13623 300
rect 13651 272 22437 300
rect 22465 272 22499 300
rect 22527 272 22561 300
rect 22589 272 22623 300
rect 22651 272 31437 300
rect 31465 272 31499 300
rect 31527 272 31561 300
rect 31589 272 31623 300
rect 31651 272 40437 300
rect 40465 272 40499 300
rect 40527 272 40561 300
rect 40589 272 40623 300
rect 40651 272 49437 300
rect 49465 272 49499 300
rect 49527 272 49561 300
rect 49589 272 49623 300
rect 49651 272 58437 300
rect 58465 272 58499 300
rect 58527 272 58561 300
rect 58589 272 58623 300
rect 58651 272 67437 300
rect 67465 272 67499 300
rect 67527 272 67561 300
rect 67589 272 67623 300
rect 67651 272 76437 300
rect 76465 272 76499 300
rect 76527 272 76561 300
rect 76589 272 76623 300
rect 76651 272 85437 300
rect 85465 272 85499 300
rect 85527 272 85561 300
rect 85589 272 85623 300
rect 85651 272 94437 300
rect 94465 272 94499 300
rect 94527 272 94561 300
rect 94589 272 94623 300
rect 94651 272 103437 300
rect 103465 272 103499 300
rect 103527 272 103561 300
rect 103589 272 103623 300
rect 103651 272 112437 300
rect 112465 272 112499 300
rect 112527 272 112561 300
rect 112589 272 112623 300
rect 112651 272 121437 300
rect 121465 272 121499 300
rect 121527 272 121561 300
rect 121589 272 121623 300
rect 121651 272 130437 300
rect 130465 272 130499 300
rect 130527 272 130561 300
rect 130589 272 130623 300
rect 130651 272 139437 300
rect 139465 272 139499 300
rect 139527 272 139561 300
rect 139589 272 139623 300
rect 139651 272 148437 300
rect 148465 272 148499 300
rect 148527 272 148561 300
rect 148589 272 148623 300
rect 148651 272 157437 300
rect 157465 272 157499 300
rect 157527 272 157561 300
rect 157589 272 157623 300
rect 157651 272 166437 300
rect 166465 272 166499 300
rect 166527 272 166561 300
rect 166589 272 166623 300
rect 166651 272 175437 300
rect 175465 272 175499 300
rect 175527 272 175561 300
rect 175589 272 175623 300
rect 175651 272 184437 300
rect 184465 272 184499 300
rect 184527 272 184561 300
rect 184589 272 184623 300
rect 184651 272 193437 300
rect 193465 272 193499 300
rect 193527 272 193561 300
rect 193589 272 193623 300
rect 193651 272 202437 300
rect 202465 272 202499 300
rect 202527 272 202561 300
rect 202589 272 202623 300
rect 202651 272 211437 300
rect 211465 272 211499 300
rect 211527 272 211561 300
rect 211589 272 211623 300
rect 211651 272 220437 300
rect 220465 272 220499 300
rect 220527 272 220561 300
rect 220589 272 220623 300
rect 220651 272 229437 300
rect 229465 272 229499 300
rect 229527 272 229561 300
rect 229589 272 229623 300
rect 229651 272 238437 300
rect 238465 272 238499 300
rect 238527 272 238561 300
rect 238589 272 238623 300
rect 238651 272 247437 300
rect 247465 272 247499 300
rect 247527 272 247561 300
rect 247589 272 247623 300
rect 247651 272 256437 300
rect 256465 272 256499 300
rect 256527 272 256561 300
rect 256589 272 256623 300
rect 256651 272 265437 300
rect 265465 272 265499 300
rect 265527 272 265561 300
rect 265589 272 265623 300
rect 265651 272 274437 300
rect 274465 272 274499 300
rect 274527 272 274561 300
rect 274589 272 274623 300
rect 274651 272 283437 300
rect 283465 272 283499 300
rect 283527 272 283561 300
rect 283589 272 283623 300
rect 283651 272 292437 300
rect 292465 272 292499 300
rect 292527 272 292561 300
rect 292589 272 292623 300
rect 292651 272 299736 300
rect 299764 272 299798 300
rect 299826 272 299860 300
rect 299888 272 299922 300
rect 299950 272 299998 300
rect -6 238 299998 272
rect -6 210 42 238
rect 70 210 104 238
rect 132 210 166 238
rect 194 210 228 238
rect 256 210 4437 238
rect 4465 210 4499 238
rect 4527 210 4561 238
rect 4589 210 4623 238
rect 4651 210 13437 238
rect 13465 210 13499 238
rect 13527 210 13561 238
rect 13589 210 13623 238
rect 13651 210 22437 238
rect 22465 210 22499 238
rect 22527 210 22561 238
rect 22589 210 22623 238
rect 22651 210 31437 238
rect 31465 210 31499 238
rect 31527 210 31561 238
rect 31589 210 31623 238
rect 31651 210 40437 238
rect 40465 210 40499 238
rect 40527 210 40561 238
rect 40589 210 40623 238
rect 40651 210 49437 238
rect 49465 210 49499 238
rect 49527 210 49561 238
rect 49589 210 49623 238
rect 49651 210 58437 238
rect 58465 210 58499 238
rect 58527 210 58561 238
rect 58589 210 58623 238
rect 58651 210 67437 238
rect 67465 210 67499 238
rect 67527 210 67561 238
rect 67589 210 67623 238
rect 67651 210 76437 238
rect 76465 210 76499 238
rect 76527 210 76561 238
rect 76589 210 76623 238
rect 76651 210 85437 238
rect 85465 210 85499 238
rect 85527 210 85561 238
rect 85589 210 85623 238
rect 85651 210 94437 238
rect 94465 210 94499 238
rect 94527 210 94561 238
rect 94589 210 94623 238
rect 94651 210 103437 238
rect 103465 210 103499 238
rect 103527 210 103561 238
rect 103589 210 103623 238
rect 103651 210 112437 238
rect 112465 210 112499 238
rect 112527 210 112561 238
rect 112589 210 112623 238
rect 112651 210 121437 238
rect 121465 210 121499 238
rect 121527 210 121561 238
rect 121589 210 121623 238
rect 121651 210 130437 238
rect 130465 210 130499 238
rect 130527 210 130561 238
rect 130589 210 130623 238
rect 130651 210 139437 238
rect 139465 210 139499 238
rect 139527 210 139561 238
rect 139589 210 139623 238
rect 139651 210 148437 238
rect 148465 210 148499 238
rect 148527 210 148561 238
rect 148589 210 148623 238
rect 148651 210 157437 238
rect 157465 210 157499 238
rect 157527 210 157561 238
rect 157589 210 157623 238
rect 157651 210 166437 238
rect 166465 210 166499 238
rect 166527 210 166561 238
rect 166589 210 166623 238
rect 166651 210 175437 238
rect 175465 210 175499 238
rect 175527 210 175561 238
rect 175589 210 175623 238
rect 175651 210 184437 238
rect 184465 210 184499 238
rect 184527 210 184561 238
rect 184589 210 184623 238
rect 184651 210 193437 238
rect 193465 210 193499 238
rect 193527 210 193561 238
rect 193589 210 193623 238
rect 193651 210 202437 238
rect 202465 210 202499 238
rect 202527 210 202561 238
rect 202589 210 202623 238
rect 202651 210 211437 238
rect 211465 210 211499 238
rect 211527 210 211561 238
rect 211589 210 211623 238
rect 211651 210 220437 238
rect 220465 210 220499 238
rect 220527 210 220561 238
rect 220589 210 220623 238
rect 220651 210 229437 238
rect 229465 210 229499 238
rect 229527 210 229561 238
rect 229589 210 229623 238
rect 229651 210 238437 238
rect 238465 210 238499 238
rect 238527 210 238561 238
rect 238589 210 238623 238
rect 238651 210 247437 238
rect 247465 210 247499 238
rect 247527 210 247561 238
rect 247589 210 247623 238
rect 247651 210 256437 238
rect 256465 210 256499 238
rect 256527 210 256561 238
rect 256589 210 256623 238
rect 256651 210 265437 238
rect 265465 210 265499 238
rect 265527 210 265561 238
rect 265589 210 265623 238
rect 265651 210 274437 238
rect 274465 210 274499 238
rect 274527 210 274561 238
rect 274589 210 274623 238
rect 274651 210 283437 238
rect 283465 210 283499 238
rect 283527 210 283561 238
rect 283589 210 283623 238
rect 283651 210 292437 238
rect 292465 210 292499 238
rect 292527 210 292561 238
rect 292589 210 292623 238
rect 292651 210 299736 238
rect 299764 210 299798 238
rect 299826 210 299860 238
rect 299888 210 299922 238
rect 299950 210 299998 238
rect -6 162 299998 210
use wrapped_rc4  rc4_1
timestamp 0
transform 1 0 15000 0 1 15000
box -28 -28 239988 239988
<< labels >>
flabel metal3 s 299760 3332 300480 3444 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 299760 203252 300480 203364 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 299760 223244 300480 223356 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 299760 243236 300480 243348 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 299760 263228 300480 263340 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 299760 283220 300480 283332 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 294084 299760 294196 300480 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 260820 299760 260932 300480 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 227556 299760 227668 300480 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 194292 299760 194404 300480 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 161028 299760 161140 300480 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 299760 23324 300480 23436 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 127764 299760 127876 300480 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 94500 299760 94612 300480 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 61236 299760 61348 300480 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 27972 299760 28084 300480 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -480 295708 240 295820 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -480 274372 240 274484 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -480 253036 240 253148 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -480 231700 240 231812 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -480 210364 240 210476 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -480 189028 240 189140 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 299760 43316 300480 43428 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -480 167692 240 167804 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -480 146356 240 146468 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -480 125020 240 125132 0 FreeSans 448 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -480 103684 240 103796 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -480 82348 240 82460 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -480 61012 240 61124 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -480 39676 240 39788 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -480 18340 240 18452 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 299760 63308 300480 63420 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 299760 83300 300480 83412 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 299760 103292 300480 103404 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 299760 123284 300480 123396 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 299760 143276 300480 143388 0 FreeSans 448 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 299760 163268 300480 163380 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 299760 183260 300480 183372 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 299760 16660 300480 16772 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 299760 216580 300480 216692 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 299760 236572 300480 236684 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 299760 256564 300480 256676 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 299760 276556 300480 276668 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 299760 296548 300480 296660 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 271908 299760 272020 300480 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 238644 299760 238756 300480 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 205380 299760 205492 300480 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 172116 299760 172228 300480 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 138852 299760 138964 300480 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 299760 36652 300480 36764 0 FreeSans 448 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 105588 299760 105700 300480 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 72324 299760 72436 300480 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 39060 299760 39172 300480 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 5796 299760 5908 300480 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -480 281484 240 281596 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -480 260148 240 260260 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -480 238812 240 238924 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -480 217476 240 217588 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -480 196140 240 196252 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -480 174804 240 174916 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 299760 56644 300480 56756 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -480 153468 240 153580 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -480 132132 240 132244 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -480 110796 240 110908 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -480 89460 240 89572 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -480 68124 240 68236 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -480 46788 240 46900 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -480 25452 240 25564 0 FreeSans 448 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -480 4116 240 4228 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 299760 76636 300480 76748 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 299760 96628 300480 96740 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 299760 116620 300480 116732 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 299760 136612 300480 136724 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 299760 156604 300480 156716 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 299760 176596 300480 176708 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 299760 196588 300480 196700 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 299760 9996 300480 10108 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 299760 209916 300480 210028 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 299760 229908 300480 230020 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 299760 249900 300480 250012 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 299760 269892 300480 270004 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 299760 289884 300480 289996 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 282996 299760 283108 300480 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 249732 299760 249844 300480 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 216468 299760 216580 300480 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 183204 299760 183316 300480 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 149940 299760 150052 300480 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 299760 29988 300480 30100 0 FreeSans 448 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 116676 299760 116788 300480 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 83412 299760 83524 300480 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 50148 299760 50260 300480 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 16884 299760 16996 300480 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -480 288596 240 288708 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -480 267260 240 267372 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -480 245924 240 246036 0 FreeSans 448 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -480 224588 240 224700 0 FreeSans 448 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -480 203252 240 203364 0 FreeSans 448 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -480 181916 240 182028 0 FreeSans 448 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 299760 49980 300480 50092 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -480 160580 240 160692 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -480 139244 240 139356 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -480 117908 240 118020 0 FreeSans 448 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -480 96572 240 96684 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -480 75236 240 75348 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -480 53900 240 54012 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -480 32564 240 32676 0 FreeSans 448 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -480 11228 240 11340 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 299760 69972 300480 70084 0 FreeSans 448 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 299760 89964 300480 90076 0 FreeSans 448 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 299760 109956 300480 110068 0 FreeSans 448 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 299760 129948 300480 130060 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 299760 149940 300480 150052 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 299760 169932 300480 170044 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 299760 189924 300480 190036 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 107548 -480 107660 240 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 136108 -480 136220 240 0 FreeSans 448 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 138964 -480 139076 240 0 FreeSans 448 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 141820 -480 141932 240 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 144676 -480 144788 240 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 147532 -480 147644 240 0 FreeSans 448 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 150388 -480 150500 240 0 FreeSans 448 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 153244 -480 153356 240 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 156100 -480 156212 240 0 FreeSans 448 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 158956 -480 159068 240 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 161812 -480 161924 240 0 FreeSans 448 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 110404 -480 110516 240 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 164668 -480 164780 240 0 FreeSans 448 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 167524 -480 167636 240 0 FreeSans 448 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 170380 -480 170492 240 0 FreeSans 448 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 173236 -480 173348 240 0 FreeSans 448 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 176092 -480 176204 240 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 178948 -480 179060 240 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 181804 -480 181916 240 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 184660 -480 184772 240 0 FreeSans 448 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 187516 -480 187628 240 0 FreeSans 448 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 190372 -480 190484 240 0 FreeSans 448 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 113260 -480 113372 240 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 193228 -480 193340 240 0 FreeSans 448 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 196084 -480 196196 240 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 198940 -480 199052 240 0 FreeSans 448 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 201796 -480 201908 240 0 FreeSans 448 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 204652 -480 204764 240 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 207508 -480 207620 240 0 FreeSans 448 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 210364 -480 210476 240 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 213220 -480 213332 240 0 FreeSans 448 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 216076 -480 216188 240 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 218932 -480 219044 240 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 116116 -480 116228 240 0 FreeSans 448 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 221788 -480 221900 240 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 224644 -480 224756 240 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 227500 -480 227612 240 0 FreeSans 448 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 230356 -480 230468 240 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 233212 -480 233324 240 0 FreeSans 448 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 236068 -480 236180 240 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 238924 -480 239036 240 0 FreeSans 448 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 241780 -480 241892 240 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 244636 -480 244748 240 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 247492 -480 247604 240 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 118972 -480 119084 240 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 250348 -480 250460 240 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 253204 -480 253316 240 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 256060 -480 256172 240 0 FreeSans 448 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 258916 -480 259028 240 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 261772 -480 261884 240 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 264628 -480 264740 240 0 FreeSans 448 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 267484 -480 267596 240 0 FreeSans 448 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 270340 -480 270452 240 0 FreeSans 448 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 273196 -480 273308 240 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 276052 -480 276164 240 0 FreeSans 448 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 121828 -480 121940 240 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 278908 -480 279020 240 0 FreeSans 448 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 281764 -480 281876 240 0 FreeSans 448 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 284620 -480 284732 240 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 287476 -480 287588 240 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 124684 -480 124796 240 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 127540 -480 127652 240 0 FreeSans 448 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 130396 -480 130508 240 0 FreeSans 448 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 133252 -480 133364 240 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 108500 -480 108612 240 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 137060 -480 137172 240 0 FreeSans 448 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 139916 -480 140028 240 0 FreeSans 448 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 142772 -480 142884 240 0 FreeSans 448 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 145628 -480 145740 240 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 148484 -480 148596 240 0 FreeSans 448 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 151340 -480 151452 240 0 FreeSans 448 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 154196 -480 154308 240 0 FreeSans 448 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 157052 -480 157164 240 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 159908 -480 160020 240 0 FreeSans 448 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 162764 -480 162876 240 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 111356 -480 111468 240 0 FreeSans 448 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 165620 -480 165732 240 0 FreeSans 448 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 168476 -480 168588 240 0 FreeSans 448 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 171332 -480 171444 240 0 FreeSans 448 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 174188 -480 174300 240 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 177044 -480 177156 240 0 FreeSans 448 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 179900 -480 180012 240 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 182756 -480 182868 240 0 FreeSans 448 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 185612 -480 185724 240 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 188468 -480 188580 240 0 FreeSans 448 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 191324 -480 191436 240 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 114212 -480 114324 240 0 FreeSans 448 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 194180 -480 194292 240 0 FreeSans 448 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 197036 -480 197148 240 0 FreeSans 448 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 199892 -480 200004 240 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 202748 -480 202860 240 0 FreeSans 448 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 205604 -480 205716 240 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 208460 -480 208572 240 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 211316 -480 211428 240 0 FreeSans 448 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 214172 -480 214284 240 0 FreeSans 448 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 217028 -480 217140 240 0 FreeSans 448 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 219884 -480 219996 240 0 FreeSans 448 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 117068 -480 117180 240 0 FreeSans 448 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 222740 -480 222852 240 0 FreeSans 448 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 225596 -480 225708 240 0 FreeSans 448 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 228452 -480 228564 240 0 FreeSans 448 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 231308 -480 231420 240 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 234164 -480 234276 240 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 237020 -480 237132 240 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 239876 -480 239988 240 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 242732 -480 242844 240 0 FreeSans 448 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 245588 -480 245700 240 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 248444 -480 248556 240 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 119924 -480 120036 240 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 251300 -480 251412 240 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 254156 -480 254268 240 0 FreeSans 448 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 257012 -480 257124 240 0 FreeSans 448 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 259868 -480 259980 240 0 FreeSans 448 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 262724 -480 262836 240 0 FreeSans 448 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 265580 -480 265692 240 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 268436 -480 268548 240 0 FreeSans 448 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 271292 -480 271404 240 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 274148 -480 274260 240 0 FreeSans 448 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 277004 -480 277116 240 0 FreeSans 448 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 122780 -480 122892 240 0 FreeSans 448 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 279860 -480 279972 240 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 282716 -480 282828 240 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 285572 -480 285684 240 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 288428 -480 288540 240 0 FreeSans 448 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 125636 -480 125748 240 0 FreeSans 448 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 128492 -480 128604 240 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 131348 -480 131460 240 0 FreeSans 448 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 134204 -480 134316 240 0 FreeSans 448 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 109452 -480 109564 240 0 FreeSans 448 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 138012 -480 138124 240 0 FreeSans 448 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 140868 -480 140980 240 0 FreeSans 448 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 143724 -480 143836 240 0 FreeSans 448 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 146580 -480 146692 240 0 FreeSans 448 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 149436 -480 149548 240 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 152292 -480 152404 240 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 155148 -480 155260 240 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 158004 -480 158116 240 0 FreeSans 448 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 160860 -480 160972 240 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 163716 -480 163828 240 0 FreeSans 448 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 112308 -480 112420 240 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 166572 -480 166684 240 0 FreeSans 448 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 169428 -480 169540 240 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 172284 -480 172396 240 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 175140 -480 175252 240 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 177996 -480 178108 240 0 FreeSans 448 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 180852 -480 180964 240 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 183708 -480 183820 240 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 186564 -480 186676 240 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 189420 -480 189532 240 0 FreeSans 448 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 192276 -480 192388 240 0 FreeSans 448 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 115164 -480 115276 240 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 195132 -480 195244 240 0 FreeSans 448 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 197988 -480 198100 240 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 200844 -480 200956 240 0 FreeSans 448 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 203700 -480 203812 240 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 206556 -480 206668 240 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 209412 -480 209524 240 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 212268 -480 212380 240 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 215124 -480 215236 240 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 217980 -480 218092 240 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 220836 -480 220948 240 0 FreeSans 448 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 118020 -480 118132 240 0 FreeSans 448 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 223692 -480 223804 240 0 FreeSans 448 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 226548 -480 226660 240 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 229404 -480 229516 240 0 FreeSans 448 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 232260 -480 232372 240 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 235116 -480 235228 240 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 237972 -480 238084 240 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 240828 -480 240940 240 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 243684 -480 243796 240 0 FreeSans 448 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 246540 -480 246652 240 0 FreeSans 448 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 249396 -480 249508 240 0 FreeSans 448 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 120876 -480 120988 240 0 FreeSans 448 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 252252 -480 252364 240 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 255108 -480 255220 240 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 257964 -480 258076 240 0 FreeSans 448 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 260820 -480 260932 240 0 FreeSans 448 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 263676 -480 263788 240 0 FreeSans 448 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 266532 -480 266644 240 0 FreeSans 448 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 269388 -480 269500 240 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 272244 -480 272356 240 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 275100 -480 275212 240 0 FreeSans 448 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 277956 -480 278068 240 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 123732 -480 123844 240 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 280812 -480 280924 240 0 FreeSans 448 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 283668 -480 283780 240 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 286524 -480 286636 240 0 FreeSans 448 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 289380 -480 289492 240 0 FreeSans 448 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 126588 -480 126700 240 0 FreeSans 448 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 129444 -480 129556 240 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 132300 -480 132412 240 0 FreeSans 448 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 135156 -480 135268 240 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 290332 -480 290444 240 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 291284 -480 291396 240 0 FreeSans 448 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 292236 -480 292348 240 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 293188 -480 293300 240 0 FreeSans 448 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s 474 642 784 299238 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 474 642 299518 952 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 474 298928 299518 299238 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 299208 642 299518 299238 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 2529 162 2839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 11529 162 11839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 20529 162 20839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 29529 162 29839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 38529 162 38839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 38529 254075 38839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 47529 162 47839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 47529 254075 47839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 56529 162 56839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 56529 254075 56839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 65529 162 65839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 65529 254075 65839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 74529 162 74839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 74529 254075 74839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 83529 162 83839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 83529 254075 83839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 92529 162 92839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 92529 254075 92839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 101529 162 101839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 101529 254394 101839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110529 162 110839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 110529 254075 110839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 119529 162 119839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 119529 254075 119839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128529 162 128839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128529 254075 128839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 137529 162 137839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 137529 254075 137839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 146529 162 146839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 146529 254075 146839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 155529 162 155839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 155529 254394 155839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 164529 162 164839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 164529 254075 164839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 173529 162 173839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 173529 254075 173839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 182529 162 182839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 182529 254075 182839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 191529 162 191839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 191529 254075 191839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 200529 162 200839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 200529 254075 200839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 209529 162 209839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 209529 254075 209839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 218529 162 218839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 218529 254075 218839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 227529 162 227839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 227529 254075 227839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 236529 162 236839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 236529 254075 236839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 245529 162 245839 14541 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 245529 254075 245839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 254529 162 254839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 263529 162 263839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 272529 162 272839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281529 162 281839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 290529 162 290839 299718 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 2697 299998 3007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 11697 299998 12007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 20697 299998 21007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 29697 299998 30007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 38697 299998 39007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 47697 299998 48007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 56697 299998 57007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 65697 299998 66007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 74697 299998 75007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 83697 299998 84007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 92697 299998 93007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 101697 299998 102007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 110697 299998 111007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 119697 299998 120007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 128697 299998 129007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 137697 299998 138007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 146697 299998 147007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 155697 299998 156007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 164697 299998 165007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 173697 299998 174007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 182697 299998 183007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 191697 299998 192007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 200697 299998 201007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 209697 299998 210007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 218697 299998 219007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 227697 299998 228007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 236697 299998 237007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 245697 299998 246007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 254697 299998 255007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 263697 299998 264007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 272697 299998 273007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 281697 299998 282007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -6 290697 299998 291007 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -6 162 304 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 162 299998 472 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 299408 299998 299718 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 299688 162 299998 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 4389 162 4699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 13389 162 13699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 22389 162 22699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 31389 162 31699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 40389 162 40699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 40389 254394 40699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 49389 162 49699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 49389 254075 49699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 58389 162 58699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 58389 254075 58699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 67389 162 67699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 67389 254075 67699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 76389 162 76699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 76389 254075 76699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 85389 162 85699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 85389 254075 85699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 94389 162 94699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 94389 254075 94699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 103389 162 103699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 103389 254075 103699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112389 162 112699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 112389 254075 112699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 121389 162 121699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 121389 254075 121699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 130389 162 130699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 130389 254075 130699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 139389 162 139699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 139389 254075 139699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 148389 162 148699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 148389 254075 148699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 157389 162 157699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 157389 254075 157699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 166389 162 166699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 166389 254075 166699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 175389 162 175699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 175389 254075 175699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 184389 162 184699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 184389 254075 184699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193389 162 193699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193389 254075 193699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 202389 162 202699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 202389 254075 202699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 211389 162 211699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 211389 254075 211699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 220389 162 220699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 220389 254075 220699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 229389 162 229699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 229389 254075 229699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 238389 162 238699 14541 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 238389 254075 238699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 247389 162 247699 15510 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 247389 254394 247699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 256389 162 256699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 265389 162 265699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 274389 162 274699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 283389 162 283699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 292389 162 292699 299718 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 5697 299998 6007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 14697 299998 15007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 23697 299998 24007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 32697 299998 33007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 41697 299998 42007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 50697 299998 51007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 59697 299998 60007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 68697 299998 69007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 77697 299998 78007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 86697 299998 87007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 95697 299998 96007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 104697 299998 105007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 113697 299998 114007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 122697 299998 123007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 131697 299998 132007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 140697 299998 141007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 149697 299998 150007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 158697 299998 159007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 167697 299998 168007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 176697 299998 177007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 185697 299998 186007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 194697 299998 195007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 203697 299998 204007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 212697 299998 213007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 221697 299998 222007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 230697 299998 231007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 239697 299998 240007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 248697 299998 249007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 257697 299998 258007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 266697 299998 267007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 275697 299998 276007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 284697 299998 285007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -6 293697 299998 294007 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 6636 -480 6748 240 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 7588 -480 7700 240 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 8540 -480 8652 240 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 12348 -480 12460 240 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 44716 -480 44828 240 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 47572 -480 47684 240 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 50428 -480 50540 240 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 53284 -480 53396 240 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 56140 -480 56252 240 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 58996 -480 59108 240 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 61852 -480 61964 240 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 64708 -480 64820 240 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 67564 -480 67676 240 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 70420 -480 70532 240 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 16156 -480 16268 240 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 73276 -480 73388 240 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 76132 -480 76244 240 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 78988 -480 79100 240 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 81844 -480 81956 240 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 84700 -480 84812 240 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 87556 -480 87668 240 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 90412 -480 90524 240 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 93268 -480 93380 240 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 96124 -480 96236 240 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 98980 -480 99092 240 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 19964 -480 20076 240 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 101836 -480 101948 240 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 104692 -480 104804 240 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 23772 -480 23884 240 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 27580 -480 27692 240 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 30436 -480 30548 240 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 33292 -480 33404 240 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 36148 -480 36260 240 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 39004 -480 39116 240 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 41860 -480 41972 240 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 9492 -480 9604 240 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 13300 -480 13412 240 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 45668 -480 45780 240 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 48524 -480 48636 240 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 51380 -480 51492 240 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 54236 -480 54348 240 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 57092 -480 57204 240 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 59948 -480 60060 240 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 62804 -480 62916 240 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 65660 -480 65772 240 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 68516 -480 68628 240 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 71372 -480 71484 240 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 17108 -480 17220 240 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 74228 -480 74340 240 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 77084 -480 77196 240 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 79940 -480 80052 240 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 82796 -480 82908 240 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 85652 -480 85764 240 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 88508 -480 88620 240 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 91364 -480 91476 240 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 94220 -480 94332 240 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 97076 -480 97188 240 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 99932 -480 100044 240 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 20916 -480 21028 240 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 102788 -480 102900 240 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 105644 -480 105756 240 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 24724 -480 24836 240 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 28532 -480 28644 240 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 31388 -480 31500 240 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 34244 -480 34356 240 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 37100 -480 37212 240 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 39956 -480 40068 240 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 42812 -480 42924 240 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 14252 -480 14364 240 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 46620 -480 46732 240 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 49476 -480 49588 240 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 52332 -480 52444 240 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 55188 -480 55300 240 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 58044 -480 58156 240 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 60900 -480 61012 240 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 63756 -480 63868 240 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 66612 -480 66724 240 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 69468 -480 69580 240 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 72324 -480 72436 240 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 18060 -480 18172 240 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 75180 -480 75292 240 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 78036 -480 78148 240 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 80892 -480 81004 240 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 83748 -480 83860 240 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 86604 -480 86716 240 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 89460 -480 89572 240 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 92316 -480 92428 240 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 95172 -480 95284 240 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 98028 -480 98140 240 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 100884 -480 100996 240 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 21868 -480 21980 240 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 103740 -480 103852 240 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 106596 -480 106708 240 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 25676 -480 25788 240 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 29484 -480 29596 240 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 32340 -480 32452 240 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 35196 -480 35308 240 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 38052 -480 38164 240 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 40908 -480 41020 240 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 43764 -480 43876 240 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 15204 -480 15316 240 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 19012 -480 19124 240 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 22820 -480 22932 240 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 26628 -480 26740 240 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 10444 -480 10556 240 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 11396 -480 11508 240 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 254777 254945 254777 254945 0 vdd
rlabel via4 247637 14945 247637 14945 0 vss
rlabel metal3 278621 3388 278621 3388 0 io_in[0]
rlabel metal3 256809 72828 256809 72828 0 io_in[10]
rlabel metal2 39564 255619 39564 255619 0 io_in[11]
rlabel metal3 13825 147420 13825 147420 0 io_in[12]
rlabel metal3 299796 263060 299796 263060 0 io_in[13]
rlabel metal3 294000 283164 294000 283164 0 io_in[14]
rlabel metal2 294084 298781 294084 298781 0 io_in[15]
rlabel metal2 260596 299796 260596 299796 0 io_in[16]
rlabel metal2 227164 299796 227164 299796 0 io_in[17]
rlabel metal2 236628 261436 236628 261436 0 io_in[18]
rlabel metal3 13013 47908 13013 47908 0 io_in[19]
rlabel metal2 259140 126448 259140 126448 0 io_in[1]
rlabel metal2 127736 294000 127736 294000 0 io_in[20]
rlabel metal2 94612 298809 94612 298809 0 io_in[21]
rlabel metal3 14749 180684 14749 180684 0 io_in[22]
rlabel metal2 27832 299796 27832 299796 0 io_in[23]
rlabel metal3 1155 295708 1155 295708 0 io_in[24]
rlabel metal3 1995 274372 1995 274372 0 io_in[25]
rlabel metal3 15148 238077 15148 238077 0 io_in[26]
rlabel metal3 1211 231812 1211 231812 0 io_in[27]
rlabel metal3 1183 210476 1183 210476 0 io_in[28]
rlabel metal3 2023 189028 2023 189028 0 io_in[29]
rlabel metal3 299796 43064 299796 43064 0 io_in[2]
rlabel metal3 2835 167804 2835 167804 0 io_in[30]
rlabel metal3 2835 146356 2835 146356 0 io_in[31]
rlabel metal3 2716 31892 2716 31892 0 io_in[32]
rlabel metal3 15148 155589 15148 155589 0 io_in[33]
rlabel metal2 72772 14777 72772 14777 0 io_in[34]
rlabel metal3 1267 61012 1267 61012 0 io_in[35]
rlabel metal3 3472 36092 3472 36092 0 io_in[36]
rlabel metal3 196 17976 196 17976 0 io_in[37]
rlabel metal3 299796 63140 299796 63140 0 io_in[3]
rlabel metal3 294000 83244 294000 83244 0 io_in[4]
rlabel metal3 256599 147420 256599 147420 0 io_in[5]
rlabel metal3 299796 122948 299796 122948 0 io_in[6]
rlabel metal3 298781 143276 298781 143276 0 io_in[7]
rlabel metal2 155820 255703 155820 255703 0 io_in[8]
rlabel metal2 262500 219352 262500 219352 0 io_in[9]
rlabel metal3 299796 9604 299796 9604 0 io_out[0]
rlabel metal3 299796 209524 299796 209524 0 io_out[10]
rlabel metal3 14637 188748 14637 188748 0 io_out[11]
rlabel metal3 299796 249676 299796 249676 0 io_out[12]
rlabel metal3 14245 139020 14245 139020 0 io_out[13]
rlabel metal3 15148 22869 15148 22869 0 io_out[14]
rlabel metal2 282996 298809 282996 298809 0 io_out[15]
rlabel metal2 249592 299796 249592 299796 0 io_out[16]
rlabel metal2 216580 298837 216580 298837 0 io_out[17]
rlabel metal3 189420 283892 189420 283892 0 io_out[18]
rlabel metal3 14721 64428 14721 64428 0 io_out[19]
rlabel metal3 14749 106036 14749 106036 0 io_out[1]
rlabel metal3 14196 15932 14196 15932 0 io_out[20]
rlabel metal3 15932 261660 15932 261660 0 io_out[21]
rlabel metal2 50148 298809 50148 298809 0 io_out[22]
rlabel metal2 16856 294000 16856 294000 0 io_out[23]
rlabel metal3 2835 288596 2835 288596 0 io_out[24]
rlabel metal3 5880 267204 5880 267204 0 io_out[25]
rlabel metal3 196 245588 196 245588 0 io_out[26]
rlabel metal3 1211 224588 1211 224588 0 io_out[27]
rlabel metal2 213388 255640 213388 255640 0 io_out[28]
rlabel metal3 1155 182028 1155 182028 0 io_out[29]
rlabel metal2 130956 14609 130956 14609 0 io_out[2]
rlabel metal3 5880 160524 5880 160524 0 io_out[30]
rlabel metal3 3360 24332 3360 24332 0 io_out[31]
rlabel metal3 196 117740 196 117740 0 io_out[32]
rlabel metal2 13468 97132 13468 97132 0 io_out[33]
rlabel metal3 196 74984 196 74984 0 io_out[34]
rlabel metal3 15260 15316 15260 15316 0 io_out[35]
rlabel metal3 196 32228 196 32228 0 io_out[36]
rlabel metal3 196 11060 196 11060 0 io_out[37]
rlabel metal2 261660 41944 261660 41944 0 io_out[3]
rlabel metal2 14280 15988 14280 15988 0 io_out[4]
rlabel metal3 299796 109564 299796 109564 0 io_out[5]
rlabel metal3 299796 129640 299796 129640 0 io_out[6]
rlabel metal2 64428 255619 64428 255619 0 io_out[7]
rlabel metal2 180684 14609 180684 14609 0 io_out[8]
rlabel metal3 14476 252028 14476 252028 0 io_out[9]
rlabel metal3 15148 221865 15148 221865 0 wb_clk_i
rlabel metal3 132356 13860 132356 13860 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 300000 300000
<< end >>
